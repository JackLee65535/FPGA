`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/06/30 10:49:38
// Design Name: 
// Module Name: mem_4096x1024
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mem_4096x1024(
    input   sclk,
    input   rst_n,
    input   en,
    input       [11:0]  addr,
    output  reg [11:0]  data
    );
    
    reg   [11:0]  mem[4095:0];
    
    
    initial begin
    mem[0] = 0;
    mem[1] = 2;
    mem[2] = 3;
    mem[3] = 5;
    mem[4] = 6;
    mem[5] = 8;
    mem[6] = 9;
    mem[7] = 11;
    mem[8] = 13;
    mem[9] = 14;
    mem[10] = 16;
    mem[11] = 17;
    mem[12] = 19;
    mem[13] = 20;
    mem[14] = 22;
    mem[15] = 24;
    mem[16] = 25;
    mem[17] = 27;
    mem[18] = 28;
    mem[19] = 30;
    mem[20] = 31;
    mem[21] = 33;
    mem[22] = 35;
    mem[23] = 36;
    mem[24] = 38;
    mem[25] = 39;
    mem[26] = 41;
    mem[27] = 42;
    mem[28] = 44;
    mem[29] = 46;
    mem[30] = 47;
    mem[31] = 49;
    mem[32] = 50;
    mem[33] = 52;
    mem[34] = 53;
    mem[35] = 55;
    mem[36] = 57;
    mem[37] = 58;
    mem[38] = 60;
    mem[39] = 61;
    mem[40] = 63;
    mem[41] = 64;
    mem[42] = 66;
    mem[43] = 68;
    mem[44] = 69;
    mem[45] = 71;
    mem[46] = 72;
    mem[47] = 74;
    mem[48] = 75;
    mem[49] = 77;
    mem[50] = 78;
    mem[51] = 80;
    mem[52] = 82;
    mem[53] = 83;
    mem[54] = 85;
    mem[55] = 86;
    mem[56] = 88;
    mem[57] = 89;
    mem[58] = 91;
    mem[59] = 93;
    mem[60] = 94;
    mem[61] = 96;
    mem[62] = 97;
    mem[63] = 99;
    mem[64] = 100;
    mem[65] = 102;
    mem[66] = 104;
    mem[67] = 105;
    mem[68] = 107;
    mem[69] = 108;
    mem[70] = 110;
    mem[71] = 111;
    mem[72] = 113;
    mem[73] = 114;
    mem[74] = 116;
    mem[75] = 118;
    mem[76] = 119;
    mem[77] = 121;
    mem[78] = 122;
    mem[79] = 124;
    mem[80] = 125;
    mem[81] = 127;
    mem[82] = 128;
    mem[83] = 130;
    mem[84] = 132;
    mem[85] = 133;
    mem[86] = 135;
    mem[87] = 136;
    mem[88] = 138;
    mem[89] = 139;
    mem[90] = 141;
    mem[91] = 143;
    mem[92] = 144;
    mem[93] = 146;
    mem[94] = 147;
    mem[95] = 149;
    mem[96] = 150;
    mem[97] = 152;
    mem[98] = 153;
    mem[99] = 155;
    mem[100] = 157;
    mem[101] = 158;
    mem[102] = 160;
    mem[103] = 161;
    mem[104] = 163;
    mem[105] = 164;
    mem[106] = 166;
    mem[107] = 167;
    mem[108] = 169;
    mem[109] = 170;
    mem[110] = 172;
    mem[111] = 174;
    mem[112] = 175;
    mem[113] = 177;
    mem[114] = 178;
    mem[115] = 180;
    mem[116] = 181;
    mem[117] = 183;
    mem[118] = 184;
    mem[119] = 186;
    mem[120] = 187;
    mem[121] = 189;
    mem[122] = 191;
    mem[123] = 192;
    mem[124] = 194;
    mem[125] = 195;
    mem[126] = 197;
    mem[127] = 198;
    mem[128] = 200;
    mem[129] = 201;
    mem[130] = 203;
    mem[131] = 204;
    mem[132] = 206;
    mem[133] = 208;
    mem[134] = 209;
    mem[135] = 211;
    mem[136] = 212;
    mem[137] = 214;
    mem[138] = 215;
    mem[139] = 217;
    mem[140] = 218;
    mem[141] = 220;
    mem[142] = 221;
    mem[143] = 223;
    mem[144] = 224;
    mem[145] = 226;
    mem[146] = 227;
    mem[147] = 229;
    mem[148] = 231;
    mem[149] = 232;
    mem[150] = 234;
    mem[151] = 235;
    mem[152] = 237;
    mem[153] = 238;
    mem[154] = 240;
    mem[155] = 241;
    mem[156] = 243;
    mem[157] = 244;
    mem[158] = 246;
    mem[159] = 247;
    mem[160] = 249;
    mem[161] = 250;
    mem[162] = 252;
    mem[163] = 253;
    mem[164] = 255;
    mem[165] = 256;
    mem[166] = 258;
    mem[167] = 260;
    mem[168] = 261;
    mem[169] = 263;
    mem[170] = 264;
    mem[171] = 266;
    mem[172] = 267;
    mem[173] = 269;
    mem[174] = 270;
    mem[175] = 272;
    mem[176] = 273;
    mem[177] = 275;
    mem[178] = 276;
    mem[179] = 278;
    mem[180] = 279;
    mem[181] = 281;
    mem[182] = 282;
    mem[183] = 284;
    mem[184] = 285;
    mem[185] = 287;
    mem[186] = 288;
    mem[187] = 290;
    mem[188] = 291;
    mem[189] = 293;
    mem[190] = 294;
    mem[191] = 296;
    mem[192] = 297;
    mem[193] = 299;
    mem[194] = 300;
    mem[195] = 302;
    mem[196] = 303;
    mem[197] = 305;
    mem[198] = 306;
    mem[199] = 308;
    mem[200] = 309;
    mem[201] = 311;
    mem[202] = 312;
    mem[203] = 314;
    mem[204] = 315;
    mem[205] = 317;
    mem[206] = 318;
    mem[207] = 320;
    mem[208] = 321;
    mem[209] = 323;
    mem[210] = 324;
    mem[211] = 326;
    mem[212] = 327;
    mem[213] = 329;
    mem[214] = 330;
    mem[215] = 332;
    mem[216] = 333;
    mem[217] = 335;
    mem[218] = 336;
    mem[219] = 338;
    mem[220] = 339;
    mem[221] = 341;
    mem[222] = 342;
    mem[223] = 344;
    mem[224] = 345;
    mem[225] = 347;
    mem[226] = 348;
    mem[227] = 349;
    mem[228] = 351;
    mem[229] = 352;
    mem[230] = 354;
    mem[231] = 355;
    mem[232] = 357;
    mem[233] = 358;
    mem[234] = 360;
    mem[235] = 361;
    mem[236] = 363;
    mem[237] = 364;
    mem[238] = 366;
    mem[239] = 367;
    mem[240] = 369;
    mem[241] = 370;
    mem[242] = 372;
    mem[243] = 373;
    mem[244] = 374;
    mem[245] = 376;
    mem[246] = 377;
    mem[247] = 379;
    mem[248] = 380;
    mem[249] = 382;
    mem[250] = 383;
    mem[251] = 385;
    mem[252] = 386;
    mem[253] = 388;
    mem[254] = 389;
    mem[255] = 391;
    mem[256] = 392;
    mem[257] = 393;
    mem[258] = 395;
    mem[259] = 396;
    mem[260] = 398;
    mem[261] = 399;
    mem[262] = 401;
    mem[263] = 402;
    mem[264] = 404;
    mem[265] = 405;
    mem[266] = 406;
    mem[267] = 408;
    mem[268] = 409;
    mem[269] = 411;
    mem[270] = 412;
    mem[271] = 414;
    mem[272] = 415;
    mem[273] = 416;
    mem[274] = 418;
    mem[275] = 419;
    mem[276] = 421;
    mem[277] = 422;
    mem[278] = 424;
    mem[279] = 425;
    mem[280] = 427;
    mem[281] = 428;
    mem[282] = 429;
    mem[283] = 431;
    mem[284] = 432;
    mem[285] = 434;
    mem[286] = 435;
    mem[287] = 436;
    mem[288] = 438;
    mem[289] = 439;
    mem[290] = 441;
    mem[291] = 442;
    mem[292] = 444;
    mem[293] = 445;
    mem[294] = 446;
    mem[295] = 448;
    mem[296] = 449;
    mem[297] = 451;
    mem[298] = 452;
    mem[299] = 453;
    mem[300] = 455;
    mem[301] = 456;
    mem[302] = 458;
    mem[303] = 459;
    mem[304] = 461;
    mem[305] = 462;
    mem[306] = 463;
    mem[307] = 465;
    mem[308] = 466;
    mem[309] = 468;
    mem[310] = 469;
    mem[311] = 470;
    mem[312] = 472;
    mem[313] = 473;
    mem[314] = 474;
    mem[315] = 476;
    mem[316] = 477;
    mem[317] = 479;
    mem[318] = 480;
    mem[319] = 481;
    mem[320] = 483;
    mem[321] = 484;
    mem[322] = 486;
    mem[323] = 487;
    mem[324] = 488;
    mem[325] = 490;
    mem[326] = 491;
    mem[327] = 492;
    mem[328] = 494;
    mem[329] = 495;
    mem[330] = 497;
    mem[331] = 498;
    mem[332] = 499;
    mem[333] = 501;
    mem[334] = 502;
    mem[335] = 503;
    mem[336] = 505;
    mem[337] = 506;
    mem[338] = 508;
    mem[339] = 509;
    mem[340] = 510;
    mem[341] = 512;
    mem[342] = 513;
    mem[343] = 514;
    mem[344] = 516;
    mem[345] = 517;
    mem[346] = 518;
    mem[347] = 520;
    mem[348] = 521;
    mem[349] = 523;
    mem[350] = 524;
    mem[351] = 525;
    mem[352] = 527;
    mem[353] = 528;
    mem[354] = 529;
    mem[355] = 531;
    mem[356] = 532;
    mem[357] = 533;
    mem[358] = 535;
    mem[359] = 536;
    mem[360] = 537;
    mem[361] = 539;
    mem[362] = 540;
    mem[363] = 541;
    mem[364] = 543;
    mem[365] = 544;
    mem[366] = 545;
    mem[367] = 547;
    mem[368] = 548;
    mem[369] = 549;
    mem[370] = 551;
    mem[371] = 552;
    mem[372] = 553;
    mem[373] = 555;
    mem[374] = 556;
    mem[375] = 557;
    mem[376] = 559;
    mem[377] = 560;
    mem[378] = 561;
    mem[379] = 562;
    mem[380] = 564;
    mem[381] = 565;
    mem[382] = 566;
    mem[383] = 568;
    mem[384] = 569;
    mem[385] = 570;
    mem[386] = 572;
    mem[387] = 573;
    mem[388] = 574;
    mem[389] = 576;
    mem[390] = 577;
    mem[391] = 578;
    mem[392] = 579;
    mem[393] = 581;
    mem[394] = 582;
    mem[395] = 583;
    mem[396] = 585;
    mem[397] = 586;
    mem[398] = 587;
    mem[399] = 588;
    mem[400] = 590;
    mem[401] = 591;
    mem[402] = 592;
    mem[403] = 594;
    mem[404] = 595;
    mem[405] = 596;
    mem[406] = 597;
    mem[407] = 599;
    mem[408] = 600;
    mem[409] = 601;
    mem[410] = 603;
    mem[411] = 604;
    mem[412] = 605;
    mem[413] = 606;
    mem[414] = 608;
    mem[415] = 609;
    mem[416] = 610;
    mem[417] = 611;
    mem[418] = 613;
    mem[419] = 614;
    mem[420] = 615;
    mem[421] = 616;
    mem[422] = 618;
    mem[423] = 619;
    mem[424] = 620;
    mem[425] = 621;
    mem[426] = 623;
    mem[427] = 624;
    mem[428] = 625;
    mem[429] = 626;
    mem[430] = 628;
    mem[431] = 629;
    mem[432] = 630;
    mem[433] = 631;
    mem[434] = 633;
    mem[435] = 634;
    mem[436] = 635;
    mem[437] = 636;
    mem[438] = 638;
    mem[439] = 639;
    mem[440] = 640;
    mem[441] = 641;
    mem[442] = 642;
    mem[443] = 644;
    mem[444] = 645;
    mem[445] = 646;
    mem[446] = 647;
    mem[447] = 649;
    mem[448] = 650;
    mem[449] = 651;
    mem[450] = 652;
    mem[451] = 653;
    mem[452] = 655;
    mem[453] = 656;
    mem[454] = 657;
    mem[455] = 658;
    mem[456] = 659;
    mem[457] = 661;
    mem[458] = 662;
    mem[459] = 663;
    mem[460] = 664;
    mem[461] = 665;
    mem[462] = 667;
    mem[463] = 668;
    mem[464] = 669;
    mem[465] = 670;
    mem[466] = 671;
    mem[467] = 673;
    mem[468] = 674;
    mem[469] = 675;
    mem[470] = 676;
    mem[471] = 677;
    mem[472] = 678;
    mem[473] = 680;
    mem[474] = 681;
    mem[475] = 682;
    mem[476] = 683;
    mem[477] = 684;
    mem[478] = 685;
    mem[479] = 687;
    mem[480] = 688;
    mem[481] = 689;
    mem[482] = 690;
    mem[483] = 691;
    mem[484] = 692;
    mem[485] = 694;
    mem[486] = 695;
    mem[487] = 696;
    mem[488] = 697;
    mem[489] = 698;
    mem[490] = 699;
    mem[491] = 701;
    mem[492] = 702;
    mem[493] = 703;
    mem[494] = 704;
    mem[495] = 705;
    mem[496] = 706;
    mem[497] = 707;
    mem[498] = 708;
    mem[499] = 710;
    mem[500] = 711;
    mem[501] = 712;
    mem[502] = 713;
    mem[503] = 714;
    mem[504] = 715;
    mem[505] = 716;
    mem[506] = 718;
    mem[507] = 719;
    mem[508] = 720;
    mem[509] = 721;
    mem[510] = 722;
    mem[511] = 723;
    mem[512] = 724;
    mem[513] = 725;
    mem[514] = 726;
    mem[515] = 728;
    mem[516] = 729;
    mem[517] = 730;
    mem[518] = 731;
    mem[519] = 732;
    mem[520] = 733;
    mem[521] = 734;
    mem[522] = 735;
    mem[523] = 736;
    mem[524] = 737;
    mem[525] = 739;
    mem[526] = 740;
    mem[527] = 741;
    mem[528] = 742;
    mem[529] = 743;
    mem[530] = 744;
    mem[531] = 745;
    mem[532] = 746;
    mem[533] = 747;
    mem[534] = 748;
    mem[535] = 749;
    mem[536] = 750;
    mem[537] = 751;
    mem[538] = 753;
    mem[539] = 754;
    mem[540] = 755;
    mem[541] = 756;
    mem[542] = 757;
    mem[543] = 758;
    mem[544] = 759;
    mem[545] = 760;
    mem[546] = 761;
    mem[547] = 762;
    mem[548] = 763;
    mem[549] = 764;
    mem[550] = 765;
    mem[551] = 766;
    mem[552] = 767;
    mem[553] = 768;
    mem[554] = 769;
    mem[555] = 770;
    mem[556] = 771;
    mem[557] = 772;
    mem[558] = 773;
    mem[559] = 774;
    mem[560] = 776;
    mem[561] = 777;
    mem[562] = 778;
    mem[563] = 779;
    mem[564] = 780;
    mem[565] = 781;
    mem[566] = 782;
    mem[567] = 783;
    mem[568] = 784;
    mem[569] = 785;
    mem[570] = 786;
    mem[571] = 787;
    mem[572] = 788;
    mem[573] = 789;
    mem[574] = 790;
    mem[575] = 791;
    mem[576] = 792;
    mem[577] = 793;
    mem[578] = 794;
    mem[579] = 795;
    mem[580] = 796;
    mem[581] = 797;
    mem[582] = 798;
    mem[583] = 799;
    mem[584] = 800;
    mem[585] = 801;
    mem[586] = 802;
    mem[587] = 803;
    mem[588] = 804;
    mem[589] = 804;
    mem[590] = 805;
    mem[591] = 806;
    mem[592] = 807;
    mem[593] = 808;
    mem[594] = 809;
    mem[595] = 810;
    mem[596] = 811;
    mem[597] = 812;
    mem[598] = 813;
    mem[599] = 814;
    mem[600] = 815;
    mem[601] = 816;
    mem[602] = 817;
    mem[603] = 818;
    mem[604] = 819;
    mem[605] = 820;
    mem[606] = 821;
    mem[607] = 822;
    mem[608] = 823;
    mem[609] = 824;
    mem[610] = 824;
    mem[611] = 825;
    mem[612] = 826;
    mem[613] = 827;
    mem[614] = 828;
    mem[615] = 829;
    mem[616] = 830;
    mem[617] = 831;
    mem[618] = 832;
    mem[619] = 833;
    mem[620] = 834;
    mem[621] = 835;
    mem[622] = 836;
    mem[623] = 836;
    mem[624] = 837;
    mem[625] = 838;
    mem[626] = 839;
    mem[627] = 840;
    mem[628] = 841;
    mem[629] = 842;
    mem[630] = 843;
    mem[631] = 844;
    mem[632] = 845;
    mem[633] = 845;
    mem[634] = 846;
    mem[635] = 847;
    mem[636] = 848;
    mem[637] = 849;
    mem[638] = 850;
    mem[639] = 851;
    mem[640] = 852;
    mem[641] = 852;
    mem[642] = 853;
    mem[643] = 854;
    mem[644] = 855;
    mem[645] = 856;
    mem[646] = 857;
    mem[647] = 858;
    mem[648] = 858;
    mem[649] = 859;
    mem[650] = 860;
    mem[651] = 861;
    mem[652] = 862;
    mem[653] = 863;
    mem[654] = 864;
    mem[655] = 864;
    mem[656] = 865;
    mem[657] = 866;
    mem[658] = 867;
    mem[659] = 868;
    mem[660] = 869;
    mem[661] = 869;
    mem[662] = 870;
    mem[663] = 871;
    mem[664] = 872;
    mem[665] = 873;
    mem[666] = 874;
    mem[667] = 874;
    mem[668] = 875;
    mem[669] = 876;
    mem[670] = 877;
    mem[671] = 878;
    mem[672] = 878;
    mem[673] = 879;
    mem[674] = 880;
    mem[675] = 881;
    mem[676] = 882;
    mem[677] = 882;
    mem[678] = 883;
    mem[679] = 884;
    mem[680] = 885;
    mem[681] = 886;
    mem[682] = 886;
    mem[683] = 887;
    mem[684] = 888;
    mem[685] = 889;
    mem[686] = 890;
    mem[687] = 890;
    mem[688] = 891;
    mem[689] = 892;
    mem[690] = 893;
    mem[691] = 893;
    mem[692] = 894;
    mem[693] = 895;
    mem[694] = 896;
    mem[695] = 896;
    mem[696] = 897;
    mem[697] = 898;
    mem[698] = 899;
    mem[699] = 899;
    mem[700] = 900;
    mem[701] = 901;
    mem[702] = 902;
    mem[703] = 902;
    mem[704] = 903;
    mem[705] = 904;
    mem[706] = 905;
    mem[707] = 905;
    mem[708] = 906;
    mem[709] = 907;
    mem[710] = 908;
    mem[711] = 908;
    mem[712] = 909;
    mem[713] = 910;
    mem[714] = 911;
    mem[715] = 911;
    mem[716] = 912;
    mem[717] = 913;
    mem[718] = 913;
    mem[719] = 914;
    mem[720] = 915;
    mem[721] = 915;
    mem[722] = 916;
    mem[723] = 917;
    mem[724] = 918;
    mem[725] = 918;
    mem[726] = 919;
    mem[727] = 920;
    mem[728] = 920;
    mem[729] = 921;
    mem[730] = 922;
    mem[731] = 922;
    mem[732] = 923;
    mem[733] = 924;
    mem[734] = 924;
    mem[735] = 925;
    mem[736] = 926;
    mem[737] = 926;
    mem[738] = 927;
    mem[739] = 928;
    mem[740] = 928;
    mem[741] = 929;
    mem[742] = 930;
    mem[743] = 930;
    mem[744] = 931;
    mem[745] = 932;
    mem[746] = 932;
    mem[747] = 933;
    mem[748] = 934;
    mem[749] = 934;
    mem[750] = 935;
    mem[751] = 936;
    mem[752] = 936;
    mem[753] = 937;
    mem[754] = 938;
    mem[755] = 938;
    mem[756] = 939;
    mem[757] = 939;
    mem[758] = 940;
    mem[759] = 941;
    mem[760] = 941;
    mem[761] = 942;
    mem[762] = 943;
    mem[763] = 943;
    mem[764] = 944;
    mem[765] = 944;
    mem[766] = 945;
    mem[767] = 946;
    mem[768] = 946;
    mem[769] = 947;
    mem[770] = 947;
    mem[771] = 948;
    mem[772] = 949;
    mem[773] = 949;
    mem[774] = 950;
    mem[775] = 950;
    mem[776] = 951;
    mem[777] = 951;
    mem[778] = 952;
    mem[779] = 953;
    mem[780] = 953;
    mem[781] = 954;
    mem[782] = 954;
    mem[783] = 955;
    mem[784] = 955;
    mem[785] = 956;
    mem[786] = 957;
    mem[787] = 957;
    mem[788] = 958;
    mem[789] = 958;
    mem[790] = 959;
    mem[791] = 959;
    mem[792] = 960;
    mem[793] = 960;
    mem[794] = 961;
    mem[795] = 962;
    mem[796] = 962;
    mem[797] = 963;
    mem[798] = 963;
    mem[799] = 964;
    mem[800] = 964;
    mem[801] = 965;
    mem[802] = 965;
    mem[803] = 966;
    mem[804] = 966;
    mem[805] = 967;
    mem[806] = 967;
    mem[807] = 968;
    mem[808] = 968;
    mem[809] = 969;
    mem[810] = 969;
    mem[811] = 970;
    mem[812] = 970;
    mem[813] = 971;
    mem[814] = 971;
    mem[815] = 972;
    mem[816] = 972;
    mem[817] = 973;
    mem[818] = 973;
    mem[819] = 974;
    mem[820] = 974;
    mem[821] = 975;
    mem[822] = 975;
    mem[823] = 976;
    mem[824] = 976;
    mem[825] = 977;
    mem[826] = 977;
    mem[827] = 978;
    mem[828] = 978;
    mem[829] = 979;
    mem[830] = 979;
    mem[831] = 980;
    mem[832] = 980;
    mem[833] = 980;
    mem[834] = 981;
    mem[835] = 981;
    mem[836] = 982;
    mem[837] = 982;
    mem[838] = 983;
    mem[839] = 983;
    mem[840] = 984;
    mem[841] = 984;
    mem[842] = 984;
    mem[843] = 985;
    mem[844] = 985;
    mem[845] = 986;
    mem[846] = 986;
    mem[847] = 987;
    mem[848] = 987;
    mem[849] = 987;
    mem[850] = 988;
    mem[851] = 988;
    mem[852] = 989;
    mem[853] = 989;
    mem[854] = 989;
    mem[855] = 990;
    mem[856] = 990;
    mem[857] = 991;
    mem[858] = 991;
    mem[859] = 991;
    mem[860] = 992;
    mem[861] = 992;
    mem[862] = 993;
    mem[863] = 993;
    mem[864] = 993;
    mem[865] = 994;
    mem[866] = 994;
    mem[867] = 995;
    mem[868] = 995;
    mem[869] = 995;
    mem[870] = 996;
    mem[871] = 996;
    mem[872] = 996;
    mem[873] = 997;
    mem[874] = 997;
    mem[875] = 997;
    mem[876] = 998;
    mem[877] = 998;
    mem[878] = 999;
    mem[879] = 999;
    mem[880] = 999;
    mem[881] = 1000;
    mem[882] = 1000;
    mem[883] = 1000;
    mem[884] = 1001;
    mem[885] = 1001;
    mem[886] = 1001;
    mem[887] = 1002;
    mem[888] = 1002;
    mem[889] = 1002;
    mem[890] = 1003;
    mem[891] = 1003;
    mem[892] = 1003;
    mem[893] = 1003;
    mem[894] = 1004;
    mem[895] = 1004;
    mem[896] = 1004;
    mem[897] = 1005;
    mem[898] = 1005;
    mem[899] = 1005;
    mem[900] = 1006;
    mem[901] = 1006;
    mem[902] = 1006;
    mem[903] = 1006;
    mem[904] = 1007;
    mem[905] = 1007;
    mem[906] = 1007;
    mem[907] = 1008;
    mem[908] = 1008;
    mem[909] = 1008;
    mem[910] = 1008;
    mem[911] = 1009;
    mem[912] = 1009;
    mem[913] = 1009;
    mem[914] = 1010;
    mem[915] = 1010;
    mem[916] = 1010;
    mem[917] = 1010;
    mem[918] = 1011;
    mem[919] = 1011;
    mem[920] = 1011;
    mem[921] = 1011;
    mem[922] = 1012;
    mem[923] = 1012;
    mem[924] = 1012;
    mem[925] = 1012;
    mem[926] = 1013;
    mem[927] = 1013;
    mem[928] = 1013;
    mem[929] = 1013;
    mem[930] = 1013;
    mem[931] = 1014;
    mem[932] = 1014;
    mem[933] = 1014;
    mem[934] = 1014;
    mem[935] = 1015;
    mem[936] = 1015;
    mem[937] = 1015;
    mem[938] = 1015;
    mem[939] = 1015;
    mem[940] = 1016;
    mem[941] = 1016;
    mem[942] = 1016;
    mem[943] = 1016;
    mem[944] = 1016;
    mem[945] = 1017;
    mem[946] = 1017;
    mem[947] = 1017;
    mem[948] = 1017;
    mem[949] = 1017;
    mem[950] = 1017;
    mem[951] = 1018;
    mem[952] = 1018;
    mem[953] = 1018;
    mem[954] = 1018;
    mem[955] = 1018;
    mem[956] = 1018;
    mem[957] = 1019;
    mem[958] = 1019;
    mem[959] = 1019;
    mem[960] = 1019;
    mem[961] = 1019;
    mem[962] = 1019;
    mem[963] = 1020;
    mem[964] = 1020;
    mem[965] = 1020;
    mem[966] = 1020;
    mem[967] = 1020;
    mem[968] = 1020;
    mem[969] = 1020;
    mem[970] = 1021;
    mem[971] = 1021;
    mem[972] = 1021;
    mem[973] = 1021;
    mem[974] = 1021;
    mem[975] = 1021;
    mem[976] = 1021;
    mem[977] = 1021;
    mem[978] = 1021;
    mem[979] = 1022;
    mem[980] = 1022;
    mem[981] = 1022;
    mem[982] = 1022;
    mem[983] = 1022;
    mem[984] = 1022;
    mem[985] = 1022;
    mem[986] = 1022;
    mem[987] = 1022;
    mem[988] = 1022;
    mem[989] = 1023;
    mem[990] = 1023;
    mem[991] = 1023;
    mem[992] = 1023;
    mem[993] = 1023;
    mem[994] = 1023;
    mem[995] = 1023;
    mem[996] = 1023;
    mem[997] = 1023;
    mem[998] = 1023;
    mem[999] = 1023;
    mem[1000] = 1023;
    mem[1001] = 1023;
    mem[1002] = 1023;
    mem[1003] = 1023;
    mem[1004] = 1024;
    mem[1005] = 1024;
    mem[1006] = 1024;
    mem[1007] = 1024;
    mem[1008] = 1024;
    mem[1009] = 1024;
    mem[1010] = 1024;
    mem[1011] = 1024;
    mem[1012] = 1024;
    mem[1013] = 1024;
    mem[1014] = 1024;
    mem[1015] = 1024;
    mem[1016] = 1024;
    mem[1017] = 1024;
    mem[1018] = 1024;
    mem[1019] = 1024;
    mem[1020] = 1024;
    mem[1021] = 1024;
    mem[1022] = 1024;
    mem[1023] = 1024;
    mem[1024] = 1024;
    mem[1025] = 1024;
    mem[1026] = 1024;
    mem[1027] = 1024;
    mem[1028] = 1024;
    mem[1029] = 1024;
    mem[1030] = 1024;
    mem[1031] = 1024;
    mem[1032] = 1024;
    mem[1033] = 1024;
    mem[1034] = 1024;
    mem[1035] = 1024;
    mem[1036] = 1024;
    mem[1037] = 1024;
    mem[1038] = 1024;
    mem[1039] = 1024;
    mem[1040] = 1024;
    mem[1041] = 1024;
    mem[1042] = 1024;
    mem[1043] = 1024;
    mem[1044] = 1024;
    mem[1045] = 1023;
    mem[1046] = 1023;
    mem[1047] = 1023;
    mem[1048] = 1023;
    mem[1049] = 1023;
    mem[1050] = 1023;
    mem[1051] = 1023;
    mem[1052] = 1023;
    mem[1053] = 1023;
    mem[1054] = 1023;
    mem[1055] = 1023;
    mem[1056] = 1023;
    mem[1057] = 1023;
    mem[1058] = 1023;
    mem[1059] = 1023;
    mem[1060] = 1022;
    mem[1061] = 1022;
    mem[1062] = 1022;
    mem[1063] = 1022;
    mem[1064] = 1022;
    mem[1065] = 1022;
    mem[1066] = 1022;
    mem[1067] = 1022;
    mem[1068] = 1022;
    mem[1069] = 1022;
    mem[1070] = 1021;
    mem[1071] = 1021;
    mem[1072] = 1021;
    mem[1073] = 1021;
    mem[1074] = 1021;
    mem[1075] = 1021;
    mem[1076] = 1021;
    mem[1077] = 1021;
    mem[1078] = 1020;
    mem[1079] = 1020;
    mem[1080] = 1020;
    mem[1081] = 1020;
    mem[1082] = 1020;
    mem[1083] = 1020;
    mem[1084] = 1020;
    mem[1085] = 1019;
    mem[1086] = 1019;
    mem[1087] = 1019;
    mem[1088] = 1019;
    mem[1089] = 1019;
    mem[1090] = 1019;
    mem[1091] = 1019;
    mem[1092] = 1018;
    mem[1093] = 1018;
    mem[1094] = 1018;
    mem[1095] = 1018;
    mem[1096] = 1018;
    mem[1097] = 1018;
    mem[1098] = 1017;
    mem[1099] = 1017;
    mem[1100] = 1017;
    mem[1101] = 1017;
    mem[1102] = 1017;
    mem[1103] = 1016;
    mem[1104] = 1016;
    mem[1105] = 1016;
    mem[1106] = 1016;
    mem[1107] = 1016;
    mem[1108] = 1015;
    mem[1109] = 1015;
    mem[1110] = 1015;
    mem[1111] = 1015;
    mem[1112] = 1015;
    mem[1113] = 1014;
    mem[1114] = 1014;
    mem[1115] = 1014;
    mem[1116] = 1014;
    mem[1117] = 1014;
    mem[1118] = 1013;
    mem[1119] = 1013;
    mem[1120] = 1013;
    mem[1121] = 1013;
    mem[1122] = 1012;
    mem[1123] = 1012;
    mem[1124] = 1012;
    mem[1125] = 1012;
    mem[1126] = 1011;
    mem[1127] = 1011;
    mem[1128] = 1011;
    mem[1129] = 1011;
    mem[1130] = 1010;
    mem[1131] = 1010;
    mem[1132] = 1010;
    mem[1133] = 1010;
    mem[1134] = 1009;
    mem[1135] = 1009;
    mem[1136] = 1009;
    mem[1137] = 1009;
    mem[1138] = 1008;
    mem[1139] = 1008;
    mem[1140] = 1008;
    mem[1141] = 1007;
    mem[1142] = 1007;
    mem[1143] = 1007;
    mem[1144] = 1007;
    mem[1145] = 1006;
    mem[1146] = 1006;
    mem[1147] = 1006;
    mem[1148] = 1005;
    mem[1149] = 1005;
    mem[1150] = 1005;
    mem[1151] = 1005;
    mem[1152] = 1004;
    mem[1153] = 1004;
    mem[1154] = 1004;
    mem[1155] = 1003;
    mem[1156] = 1003;
    mem[1157] = 1003;
    mem[1158] = 1002;
    mem[1159] = 1002;
    mem[1160] = 1002;
    mem[1161] = 1001;
    mem[1162] = 1001;
    mem[1163] = 1001;
    mem[1164] = 1000;
    mem[1165] = 1000;
    mem[1166] = 1000;
    mem[1167] = 999;
    mem[1168] = 999;
    mem[1169] = 999;
    mem[1170] = 998;
    mem[1171] = 998;
    mem[1172] = 998;
    mem[1173] = 997;
    mem[1174] = 997;
    mem[1175] = 997;
    mem[1176] = 996;
    mem[1177] = 996;
    mem[1178] = 995;
    mem[1179] = 995;
    mem[1180] = 995;
    mem[1181] = 994;
    mem[1182] = 994;
    mem[1183] = 994;
    mem[1184] = 993;
    mem[1185] = 993;
    mem[1186] = 992;
    mem[1187] = 992;
    mem[1188] = 992;
    mem[1189] = 991;
    mem[1190] = 991;
    mem[1191] = 990;
    mem[1192] = 990;
    mem[1193] = 990;
    mem[1194] = 989;
    mem[1195] = 989;
    mem[1196] = 988;
    mem[1197] = 988;
    mem[1198] = 988;
    mem[1199] = 987;
    mem[1200] = 987;
    mem[1201] = 986;
    mem[1202] = 986;
    mem[1203] = 986;
    mem[1204] = 985;
    mem[1205] = 985;
    mem[1206] = 984;
    mem[1207] = 984;
    mem[1208] = 983;
    mem[1209] = 983;
    mem[1210] = 982;
    mem[1211] = 982;
    mem[1212] = 982;
    mem[1213] = 981;
    mem[1214] = 981;
    mem[1215] = 980;
    mem[1216] = 980;
    mem[1217] = 979;
    mem[1218] = 979;
    mem[1219] = 978;
    mem[1220] = 978;
    mem[1221] = 977;
    mem[1222] = 977;
    mem[1223] = 977;
    mem[1224] = 976;
    mem[1225] = 976;
    mem[1226] = 975;
    mem[1227] = 975;
    mem[1228] = 974;
    mem[1229] = 974;
    mem[1230] = 973;
    mem[1231] = 973;
    mem[1232] = 972;
    mem[1233] = 972;
    mem[1234] = 971;
    mem[1235] = 971;
    mem[1236] = 970;
    mem[1237] = 970;
    mem[1238] = 969;
    mem[1239] = 969;
    mem[1240] = 968;
    mem[1241] = 968;
    mem[1242] = 967;
    mem[1243] = 967;
    mem[1244] = 966;
    mem[1245] = 966;
    mem[1246] = 965;
    mem[1247] = 965;
    mem[1248] = 964;
    mem[1249] = 963;
    mem[1250] = 963;
    mem[1251] = 962;
    mem[1252] = 962;
    mem[1253] = 961;
    mem[1254] = 961;
    mem[1255] = 960;
    mem[1256] = 960;
    mem[1257] = 959;
    mem[1258] = 959;
    mem[1259] = 958;
    mem[1260] = 957;
    mem[1261] = 957;
    mem[1262] = 956;
    mem[1263] = 956;
    mem[1264] = 955;
    mem[1265] = 955;
    mem[1266] = 954;
    mem[1267] = 954;
    mem[1268] = 953;
    mem[1269] = 952;
    mem[1270] = 952;
    mem[1271] = 951;
    mem[1272] = 951;
    mem[1273] = 950;
    mem[1274] = 949;
    mem[1275] = 949;
    mem[1276] = 948;
    mem[1277] = 948;
    mem[1278] = 947;
    mem[1279] = 946;
    mem[1280] = 946;
    mem[1281] = 945;
    mem[1282] = 945;
    mem[1283] = 944;
    mem[1284] = 943;
    mem[1285] = 943;
    mem[1286] = 942;
    mem[1287] = 942;
    mem[1288] = 941;
    mem[1289] = 940;
    mem[1290] = 940;
    mem[1291] = 939;
    mem[1292] = 938;
    mem[1293] = 938;
    mem[1294] = 937;
    mem[1295] = 937;
    mem[1296] = 936;
    mem[1297] = 935;
    mem[1298] = 935;
    mem[1299] = 934;
    mem[1300] = 933;
    mem[1301] = 933;
    mem[1302] = 932;
    mem[1303] = 931;
    mem[1304] = 931;
    mem[1305] = 930;
    mem[1306] = 929;
    mem[1307] = 929;
    mem[1308] = 928;
    mem[1309] = 927;
    mem[1310] = 927;
    mem[1311] = 926;
    mem[1312] = 925;
    mem[1313] = 925;
    mem[1314] = 924;
    mem[1315] = 923;
    mem[1316] = 923;
    mem[1317] = 922;
    mem[1318] = 921;
    mem[1319] = 921;
    mem[1320] = 920;
    mem[1321] = 919;
    mem[1322] = 919;
    mem[1323] = 918;
    mem[1324] = 917;
    mem[1325] = 917;
    mem[1326] = 916;
    mem[1327] = 915;
    mem[1328] = 914;
    mem[1329] = 914;
    mem[1330] = 913;
    mem[1331] = 912;
    mem[1332] = 912;
    mem[1333] = 911;
    mem[1334] = 910;
    mem[1335] = 909;
    mem[1336] = 909;
    mem[1337] = 908;
    mem[1338] = 907;
    mem[1339] = 907;
    mem[1340] = 906;
    mem[1341] = 905;
    mem[1342] = 904;
    mem[1343] = 904;
    mem[1344] = 903;
    mem[1345] = 902;
    mem[1346] = 901;
    mem[1347] = 901;
    mem[1348] = 900;
    mem[1349] = 899;
    mem[1350] = 898;
    mem[1351] = 898;
    mem[1352] = 897;
    mem[1353] = 896;
    mem[1354] = 895;
    mem[1355] = 895;
    mem[1356] = 894;
    mem[1357] = 893;
    mem[1358] = 892;
    mem[1359] = 891;
    mem[1360] = 891;
    mem[1361] = 890;
    mem[1362] = 889;
    mem[1363] = 888;
    mem[1364] = 888;
    mem[1365] = 887;
    mem[1366] = 886;
    mem[1367] = 885;
    mem[1368] = 884;
    mem[1369] = 884;
    mem[1370] = 883;
    mem[1371] = 882;
    mem[1372] = 881;
    mem[1373] = 880;
    mem[1374] = 880;
    mem[1375] = 879;
    mem[1376] = 878;
    mem[1377] = 877;
    mem[1378] = 876;
    mem[1379] = 876;
    mem[1380] = 875;
    mem[1381] = 874;
    mem[1382] = 873;
    mem[1383] = 872;
    mem[1384] = 872;
    mem[1385] = 871;
    mem[1386] = 870;
    mem[1387] = 869;
    mem[1388] = 868;
    mem[1389] = 867;
    mem[1390] = 867;
    mem[1391] = 866;
    mem[1392] = 865;
    mem[1393] = 864;
    mem[1394] = 863;
    mem[1395] = 862;
    mem[1396] = 861;
    mem[1397] = 861;
    mem[1398] = 860;
    mem[1399] = 859;
    mem[1400] = 858;
    mem[1401] = 857;
    mem[1402] = 856;
    mem[1403] = 855;
    mem[1404] = 855;
    mem[1405] = 854;
    mem[1406] = 853;
    mem[1407] = 852;
    mem[1408] = 851;
    mem[1409] = 850;
    mem[1410] = 849;
    mem[1411] = 848;
    mem[1412] = 848;
    mem[1413] = 847;
    mem[1414] = 846;
    mem[1415] = 845;
    mem[1416] = 844;
    mem[1417] = 843;
    mem[1418] = 842;
    mem[1419] = 841;
    mem[1420] = 840;
    mem[1421] = 840;
    mem[1422] = 839;
    mem[1423] = 838;
    mem[1424] = 837;
    mem[1425] = 836;
    mem[1426] = 835;
    mem[1427] = 834;
    mem[1428] = 833;
    mem[1429] = 832;
    mem[1430] = 831;
    mem[1431] = 831;
    mem[1432] = 830;
    mem[1433] = 829;
    mem[1434] = 828;
    mem[1435] = 827;
    mem[1436] = 826;
    mem[1437] = 825;
    mem[1438] = 824;
    mem[1439] = 823;
    mem[1440] = 822;
    mem[1441] = 821;
    mem[1442] = 820;
    mem[1443] = 819;
    mem[1444] = 818;
    mem[1445] = 817;
    mem[1446] = 817;
    mem[1447] = 816;
    mem[1448] = 815;
    mem[1449] = 814;
    mem[1450] = 813;
    mem[1451] = 812;
    mem[1452] = 811;
    mem[1453] = 810;
    mem[1454] = 809;
    mem[1455] = 808;
    mem[1456] = 807;
    mem[1457] = 806;
    mem[1458] = 805;
    mem[1459] = 804;
    mem[1460] = 803;
    mem[1461] = 802;
    mem[1462] = 801;
    mem[1463] = 800;
    mem[1464] = 799;
    mem[1465] = 798;
    mem[1466] = 797;
    mem[1467] = 796;
    mem[1468] = 795;
    mem[1469] = 794;
    mem[1470] = 793;
    mem[1471] = 792;
    mem[1472] = 791;
    mem[1473] = 790;
    mem[1474] = 789;
    mem[1475] = 788;
    mem[1476] = 787;
    mem[1477] = 786;
    mem[1478] = 785;
    mem[1479] = 784;
    mem[1480] = 783;
    mem[1481] = 782;
    mem[1482] = 781;
    mem[1483] = 780;
    mem[1484] = 779;
    mem[1485] = 778;
    mem[1486] = 777;
    mem[1487] = 776;
    mem[1488] = 775;
    mem[1489] = 774;
    mem[1490] = 773;
    mem[1491] = 772;
    mem[1492] = 771;
    mem[1493] = 770;
    mem[1494] = 769;
    mem[1495] = 768;
    mem[1496] = 767;
    mem[1497] = 766;
    mem[1498] = 765;
    mem[1499] = 764;
    mem[1500] = 763;
    mem[1501] = 762;
    mem[1502] = 760;
    mem[1503] = 759;
    mem[1504] = 758;
    mem[1505] = 757;
    mem[1506] = 756;
    mem[1507] = 755;
    mem[1508] = 754;
    mem[1509] = 753;
    mem[1510] = 752;
    mem[1511] = 751;
    mem[1512] = 750;
    mem[1513] = 749;
    mem[1514] = 748;
    mem[1515] = 747;
    mem[1516] = 746;
    mem[1517] = 744;
    mem[1518] = 743;
    mem[1519] = 742;
    mem[1520] = 741;
    mem[1521] = 740;
    mem[1522] = 739;
    mem[1523] = 738;
    mem[1524] = 737;
    mem[1525] = 736;
    mem[1526] = 735;
    mem[1527] = 734;
    mem[1528] = 732;
    mem[1529] = 731;
    mem[1530] = 730;
    mem[1531] = 729;
    mem[1532] = 728;
    mem[1533] = 727;
    mem[1534] = 726;
    mem[1535] = 725;
    mem[1536] = 724;
    mem[1537] = 723;
    mem[1538] = 721;
    mem[1539] = 720;
    mem[1540] = 719;
    mem[1541] = 718;
    mem[1542] = 717;
    mem[1543] = 716;
    mem[1544] = 715;
    mem[1545] = 714;
    mem[1546] = 712;
    mem[1547] = 711;
    mem[1548] = 710;
    mem[1549] = 709;
    mem[1550] = 708;
    mem[1551] = 707;
    mem[1552] = 706;
    mem[1553] = 705;
    mem[1554] = 703;
    mem[1555] = 702;
    mem[1556] = 701;
    mem[1557] = 700;
    mem[1558] = 699;
    mem[1559] = 698;
    mem[1560] = 696;
    mem[1561] = 695;
    mem[1562] = 694;
    mem[1563] = 693;
    mem[1564] = 692;
    mem[1565] = 691;
    mem[1566] = 690;
    mem[1567] = 688;
    mem[1568] = 687;
    mem[1569] = 686;
    mem[1570] = 685;
    mem[1571] = 684;
    mem[1572] = 683;
    mem[1573] = 681;
    mem[1574] = 680;
    mem[1575] = 679;
    mem[1576] = 678;
    mem[1577] = 677;
    mem[1578] = 676;
    mem[1579] = 674;
    mem[1580] = 673;
    mem[1581] = 672;
    mem[1582] = 671;
    mem[1583] = 670;
    mem[1584] = 668;
    mem[1585] = 667;
    mem[1586] = 666;
    mem[1587] = 665;
    mem[1588] = 664;
    mem[1589] = 662;
    mem[1590] = 661;
    mem[1591] = 660;
    mem[1592] = 659;
    mem[1593] = 658;
    mem[1594] = 656;
    mem[1595] = 655;
    mem[1596] = 654;
    mem[1597] = 653;
    mem[1598] = 652;
    mem[1599] = 650;
    mem[1600] = 649;
    mem[1601] = 648;
    mem[1602] = 647;
    mem[1603] = 645;
    mem[1604] = 644;
    mem[1605] = 643;
    mem[1606] = 642;
    mem[1607] = 641;
    mem[1608] = 639;
    mem[1609] = 638;
    mem[1610] = 637;
    mem[1611] = 636;
    mem[1612] = 634;
    mem[1613] = 633;
    mem[1614] = 632;
    mem[1615] = 631;
    mem[1616] = 630;
    mem[1617] = 628;
    mem[1618] = 627;
    mem[1619] = 626;
    mem[1620] = 625;
    mem[1621] = 623;
    mem[1622] = 622;
    mem[1623] = 621;
    mem[1624] = 620;
    mem[1625] = 618;
    mem[1626] = 617;
    mem[1627] = 616;
    mem[1628] = 615;
    mem[1629] = 613;
    mem[1630] = 612;
    mem[1631] = 611;
    mem[1632] = 609;
    mem[1633] = 608;
    mem[1634] = 607;
    mem[1635] = 606;
    mem[1636] = 604;
    mem[1637] = 603;
    mem[1638] = 602;
    mem[1639] = 601;
    mem[1640] = 599;
    mem[1641] = 598;
    mem[1642] = 597;
    mem[1643] = 596;
    mem[1644] = 594;
    mem[1645] = 593;
    mem[1646] = 592;
    mem[1647] = 590;
    mem[1648] = 589;
    mem[1649] = 588;
    mem[1650] = 587;
    mem[1651] = 585;
    mem[1652] = 584;
    mem[1653] = 583;
    mem[1654] = 581;
    mem[1655] = 580;
    mem[1656] = 579;
    mem[1657] = 577;
    mem[1658] = 576;
    mem[1659] = 575;
    mem[1660] = 574;
    mem[1661] = 572;
    mem[1662] = 571;
    mem[1663] = 570;
    mem[1664] = 568;
    mem[1665] = 567;
    mem[1666] = 566;
    mem[1667] = 564;
    mem[1668] = 563;
    mem[1669] = 562;
    mem[1670] = 561;
    mem[1671] = 559;
    mem[1672] = 558;
    mem[1673] = 557;
    mem[1674] = 555;
    mem[1675] = 554;
    mem[1676] = 553;
    mem[1677] = 551;
    mem[1678] = 550;
    mem[1679] = 549;
    mem[1680] = 547;
    mem[1681] = 546;
    mem[1682] = 545;
    mem[1683] = 543;
    mem[1684] = 542;
    mem[1685] = 541;
    mem[1686] = 539;
    mem[1687] = 538;
    mem[1688] = 537;
    mem[1689] = 535;
    mem[1690] = 534;
    mem[1691] = 533;
    mem[1692] = 531;
    mem[1693] = 530;
    mem[1694] = 529;
    mem[1695] = 527;
    mem[1696] = 526;
    mem[1697] = 525;
    mem[1698] = 523;
    mem[1699] = 522;
    mem[1700] = 520;
    mem[1701] = 519;
    mem[1702] = 518;
    mem[1703] = 516;
    mem[1704] = 515;
    mem[1705] = 514;
    mem[1706] = 512;
    mem[1707] = 511;
    mem[1708] = 510;
    mem[1709] = 508;
    mem[1710] = 507;
    mem[1711] = 506;
    mem[1712] = 504;
    mem[1713] = 503;
    mem[1714] = 501;
    mem[1715] = 500;
    mem[1716] = 499;
    mem[1717] = 497;
    mem[1718] = 496;
    mem[1719] = 495;
    mem[1720] = 493;
    mem[1721] = 492;
    mem[1722] = 490;
    mem[1723] = 489;
    mem[1724] = 488;
    mem[1725] = 486;
    mem[1726] = 485;
    mem[1727] = 484;
    mem[1728] = 482;
    mem[1729] = 481;
    mem[1730] = 479;
    mem[1731] = 478;
    mem[1732] = 477;
    mem[1733] = 475;
    mem[1734] = 474;
    mem[1735] = 472;
    mem[1736] = 471;
    mem[1737] = 470;
    mem[1738] = 468;
    mem[1739] = 467;
    mem[1740] = 465;
    mem[1741] = 464;
    mem[1742] = 463;
    mem[1743] = 461;
    mem[1744] = 460;
    mem[1745] = 458;
    mem[1746] = 457;
    mem[1747] = 456;
    mem[1748] = 454;
    mem[1749] = 453;
    mem[1750] = 451;
    mem[1751] = 450;
    mem[1752] = 449;
    mem[1753] = 447;
    mem[1754] = 446;
    mem[1755] = 444;
    mem[1756] = 443;
    mem[1757] = 441;
    mem[1758] = 440;
    mem[1759] = 439;
    mem[1760] = 437;
    mem[1761] = 436;
    mem[1762] = 434;
    mem[1763] = 433;
    mem[1764] = 432;
    mem[1765] = 430;
    mem[1766] = 429;
    mem[1767] = 427;
    mem[1768] = 426;
    mem[1769] = 424;
    mem[1770] = 423;
    mem[1771] = 422;
    mem[1772] = 420;
    mem[1773] = 419;
    mem[1774] = 417;
    mem[1775] = 416;
    mem[1776] = 414;
    mem[1777] = 413;
    mem[1778] = 411;
    mem[1779] = 410;
    mem[1780] = 409;
    mem[1781] = 407;
    mem[1782] = 406;
    mem[1783] = 404;
    mem[1784] = 403;
    mem[1785] = 401;
    mem[1786] = 400;
    mem[1787] = 398;
    mem[1788] = 397;
    mem[1789] = 396;
    mem[1790] = 394;
    mem[1791] = 393;
    mem[1792] = 391;
    mem[1793] = 390;
    mem[1794] = 388;
    mem[1795] = 387;
    mem[1796] = 385;
    mem[1797] = 384;
    mem[1798] = 383;
    mem[1799] = 381;
    mem[1800] = 380;
    mem[1801] = 378;
    mem[1802] = 377;
    mem[1803] = 375;
    mem[1804] = 374;
    mem[1805] = 372;
    mem[1806] = 371;
    mem[1807] = 369;
    mem[1808] = 368;
    mem[1809] = 366;
    mem[1810] = 365;
    mem[1811] = 363;
    mem[1812] = 362;
    mem[1813] = 361;
    mem[1814] = 359;
    mem[1815] = 358;
    mem[1816] = 356;
    mem[1817] = 355;
    mem[1818] = 353;
    mem[1819] = 352;
    mem[1820] = 350;
    mem[1821] = 349;
    mem[1822] = 347;
    mem[1823] = 346;
    mem[1824] = 344;
    mem[1825] = 343;
    mem[1826] = 341;
    mem[1827] = 340;
    mem[1828] = 338;
    mem[1829] = 337;
    mem[1830] = 335;
    mem[1831] = 334;
    mem[1832] = 332;
    mem[1833] = 331;
    mem[1834] = 329;
    mem[1835] = 328;
    mem[1836] = 327;
    mem[1837] = 325;
    mem[1838] = 324;
    mem[1839] = 322;
    mem[1840] = 321;
    mem[1841] = 319;
    mem[1842] = 318;
    mem[1843] = 316;
    mem[1844] = 315;
    mem[1845] = 313;
    mem[1846] = 312;
    mem[1847] = 310;
    mem[1848] = 309;
    mem[1849] = 307;
    mem[1850] = 306;
    mem[1851] = 304;
    mem[1852] = 303;
    mem[1853] = 301;
    mem[1854] = 300;
    mem[1855] = 298;
    mem[1856] = 297;
    mem[1857] = 295;
    mem[1858] = 294;
    mem[1859] = 292;
    mem[1860] = 291;
    mem[1861] = 289;
    mem[1862] = 288;
    mem[1863] = 286;
    mem[1864] = 285;
    mem[1865] = 283;
    mem[1866] = 281;
    mem[1867] = 280;
    mem[1868] = 278;
    mem[1869] = 277;
    mem[1870] = 275;
    mem[1871] = 274;
    mem[1872] = 272;
    mem[1873] = 271;
    mem[1874] = 269;
    mem[1875] = 268;
    mem[1876] = 266;
    mem[1877] = 265;
    mem[1878] = 263;
    mem[1879] = 262;
    mem[1880] = 260;
    mem[1881] = 259;
    mem[1882] = 257;
    mem[1883] = 256;
    mem[1884] = 254;
    mem[1885] = 253;
    mem[1886] = 251;
    mem[1887] = 250;
    mem[1888] = 248;
    mem[1889] = 247;
    mem[1890] = 245;
    mem[1891] = 244;
    mem[1892] = 242;
    mem[1893] = 240;
    mem[1894] = 239;
    mem[1895] = 237;
    mem[1896] = 236;
    mem[1897] = 234;
    mem[1898] = 233;
    mem[1899] = 231;
    mem[1900] = 230;
    mem[1901] = 228;
    mem[1902] = 227;
    mem[1903] = 225;
    mem[1904] = 224;
    mem[1905] = 222;
    mem[1906] = 221;
    mem[1907] = 219;
    mem[1908] = 218;
    mem[1909] = 216;
    mem[1910] = 214;
    mem[1911] = 213;
    mem[1912] = 211;
    mem[1913] = 210;
    mem[1914] = 208;
    mem[1915] = 207;
    mem[1916] = 205;
    mem[1917] = 204;
    mem[1918] = 202;
    mem[1919] = 201;
    mem[1920] = 199;
    mem[1921] = 198;
    mem[1922] = 196;
    mem[1923] = 194;
    mem[1924] = 193;
    mem[1925] = 191;
    mem[1926] = 190;
    mem[1927] = 188;
    mem[1928] = 187;
    mem[1929] = 185;
    mem[1930] = 184;
    mem[1931] = 182;
    mem[1932] = 181;
    mem[1933] = 179;
    mem[1934] = 177;
    mem[1935] = 176;
    mem[1936] = 174;
    mem[1937] = 173;
    mem[1938] = 171;
    mem[1939] = 170;
    mem[1940] = 168;
    mem[1941] = 167;
    mem[1942] = 165;
    mem[1943] = 163;
    mem[1944] = 162;
    mem[1945] = 160;
    mem[1946] = 159;
    mem[1947] = 157;
    mem[1948] = 156;
    mem[1949] = 154;
    mem[1950] = 153;
    mem[1951] = 151;
    mem[1952] = 150;
    mem[1953] = 148;
    mem[1954] = 146;
    mem[1955] = 145;
    mem[1956] = 143;
    mem[1957] = 142;
    mem[1958] = 140;
    mem[1959] = 139;
    mem[1960] = 137;
    mem[1961] = 136;
    mem[1962] = 134;
    mem[1963] = 132;
    mem[1964] = 131;
    mem[1965] = 129;
    mem[1966] = 128;
    mem[1967] = 126;
    mem[1968] = 125;
    mem[1969] = 123;
    mem[1970] = 121;
    mem[1971] = 120;
    mem[1972] = 118;
    mem[1973] = 117;
    mem[1974] = 115;
    mem[1975] = 114;
    mem[1976] = 112;
    mem[1977] = 111;
    mem[1978] = 109;
    mem[1979] = 107;
    mem[1980] = 106;
    mem[1981] = 104;
    mem[1982] = 103;
    mem[1983] = 101;
    mem[1984] = 100;
    mem[1985] = 98;
    mem[1986] = 96;
    mem[1987] = 95;
    mem[1988] = 93;
    mem[1989] = 92;
    mem[1990] = 90;
    mem[1991] = 89;
    mem[1992] = 87;
    mem[1993] = 86;
    mem[1994] = 84;
    mem[1995] = 82;
    mem[1996] = 81;
    mem[1997] = 79;
    mem[1998] = 78;
    mem[1999] = 76;
    mem[2000] = 75;
    mem[2001] = 73;
    mem[2002] = 71;
    mem[2003] = 70;
    mem[2004] = 68;
    mem[2005] = 67;
    mem[2006] = 65;
    mem[2007] = 64;
    mem[2008] = 62;
    mem[2009] = 60;
    mem[2010] = 59;
    mem[2011] = 57;
    mem[2012] = 56;
    mem[2013] = 54;
    mem[2014] = 53;
    mem[2015] = 51;
    mem[2016] = 49;
    mem[2017] = 48;
    mem[2018] = 46;
    mem[2019] = 45;
    mem[2020] = 43;
    mem[2021] = 42;
    mem[2022] = 40;
    mem[2023] = 38;
    mem[2024] = 37;
    mem[2025] = 35;
    mem[2026] = 34;
    mem[2027] = 32;
    mem[2028] = 31;
    mem[2029] = 29;
    mem[2030] = 27;
    mem[2031] = 26;
    mem[2032] = 24;
    mem[2033] = 23;
    mem[2034] = 21;
    mem[2035] = 20;
    mem[2036] = 18;
    mem[2037] = 16;
    mem[2038] = 15;
    mem[2039] = 13;
    mem[2040] = 12;
    mem[2041] = 10;
    mem[2042] = 9;
    mem[2043] = 7;
    mem[2044] = 5;
    mem[2045] = 4;
    mem[2046] = 2;
    mem[2047] = 1;
    mem[2048] = -1;
    mem[2049] = -2;
    mem[2050] = -4;
    mem[2051] = -5;
    mem[2052] = -7;
    mem[2053] = -9;
    mem[2054] = -10;
    mem[2055] = -12;
    mem[2056] = -13;
    mem[2057] = -15;
    mem[2058] = -16;
    mem[2059] = -18;
    mem[2060] = -20;
    mem[2061] = -21;
    mem[2062] = -23;
    mem[2063] = -24;
    mem[2064] = -26;
    mem[2065] = -27;
    mem[2066] = -29;
    mem[2067] = -31;
    mem[2068] = -32;
    mem[2069] = -34;
    mem[2070] = -35;
    mem[2071] = -37;
    mem[2072] = -38;
    mem[2073] = -40;
    mem[2074] = -42;
    mem[2075] = -43;
    mem[2076] = -45;
    mem[2077] = -46;
    mem[2078] = -48;
    mem[2079] = -49;
    mem[2080] = -51;
    mem[2081] = -53;
    mem[2082] = -54;
    mem[2083] = -56;
    mem[2084] = -57;
    mem[2085] = -59;
    mem[2086] = -60;
    mem[2087] = -62;
    mem[2088] = -64;
    mem[2089] = -65;
    mem[2090] = -67;
    mem[2091] = -68;
    mem[2092] = -70;
    mem[2093] = -71;
    mem[2094] = -73;
    mem[2095] = -75;
    mem[2096] = -76;
    mem[2097] = -78;
    mem[2098] = -79;
    mem[2099] = -81;
    mem[2100] = -82;
    mem[2101] = -84;
    mem[2102] = -86;
    mem[2103] = -87;
    mem[2104] = -89;
    mem[2105] = -90;
    mem[2106] = -92;
    mem[2107] = -93;
    mem[2108] = -95;
    mem[2109] = -96;
    mem[2110] = -98;
    mem[2111] = -100;
    mem[2112] = -101;
    mem[2113] = -103;
    mem[2114] = -104;
    mem[2115] = -106;
    mem[2116] = -107;
    mem[2117] = -109;
    mem[2118] = -111;
    mem[2119] = -112;
    mem[2120] = -114;
    mem[2121] = -115;
    mem[2122] = -117;
    mem[2123] = -118;
    mem[2124] = -120;
    mem[2125] = -121;
    mem[2126] = -123;
    mem[2127] = -125;
    mem[2128] = -126;
    mem[2129] = -128;
    mem[2130] = -129;
    mem[2131] = -131;
    mem[2132] = -132;
    mem[2133] = -134;
    mem[2134] = -136;
    mem[2135] = -137;
    mem[2136] = -139;
    mem[2137] = -140;
    mem[2138] = -142;
    mem[2139] = -143;
    mem[2140] = -145;
    mem[2141] = -146;
    mem[2142] = -148;
    mem[2143] = -150;
    mem[2144] = -151;
    mem[2145] = -153;
    mem[2146] = -154;
    mem[2147] = -156;
    mem[2148] = -157;
    mem[2149] = -159;
    mem[2150] = -160;
    mem[2151] = -162;
    mem[2152] = -163;
    mem[2153] = -165;
    mem[2154] = -167;
    mem[2155] = -168;
    mem[2156] = -170;
    mem[2157] = -171;
    mem[2158] = -173;
    mem[2159] = -174;
    mem[2160] = -176;
    mem[2161] = -177;
    mem[2162] = -179;
    mem[2163] = -181;
    mem[2164] = -182;
    mem[2165] = -184;
    mem[2166] = -185;
    mem[2167] = -187;
    mem[2168] = -188;
    mem[2169] = -190;
    mem[2170] = -191;
    mem[2171] = -193;
    mem[2172] = -194;
    mem[2173] = -196;
    mem[2174] = -198;
    mem[2175] = -199;
    mem[2176] = -201;
    mem[2177] = -202;
    mem[2178] = -204;
    mem[2179] = -205;
    mem[2180] = -207;
    mem[2181] = -208;
    mem[2182] = -210;
    mem[2183] = -211;
    mem[2184] = -213;
    mem[2185] = -214;
    mem[2186] = -216;
    mem[2187] = -218;
    mem[2188] = -219;
    mem[2189] = -221;
    mem[2190] = -222;
    mem[2191] = -224;
    mem[2192] = -225;
    mem[2193] = -227;
    mem[2194] = -228;
    mem[2195] = -230;
    mem[2196] = -231;
    mem[2197] = -233;
    mem[2198] = -234;
    mem[2199] = -236;
    mem[2200] = -237;
    mem[2201] = -239;
    mem[2202] = -240;
    mem[2203] = -242;
    mem[2204] = -244;
    mem[2205] = -245;
    mem[2206] = -247;
    mem[2207] = -248;
    mem[2208] = -250;
    mem[2209] = -251;
    mem[2210] = -253;
    mem[2211] = -254;
    mem[2212] = -256;
    mem[2213] = -257;
    mem[2214] = -259;
    mem[2215] = -260;
    mem[2216] = -262;
    mem[2217] = -263;
    mem[2218] = -265;
    mem[2219] = -266;
    mem[2220] = -268;
    mem[2221] = -269;
    mem[2222] = -271;
    mem[2223] = -272;
    mem[2224] = -274;
    mem[2225] = -275;
    mem[2226] = -277;
    mem[2227] = -278;
    mem[2228] = -280;
    mem[2229] = -281;
    mem[2230] = -283;
    mem[2231] = -285;
    mem[2232] = -286;
    mem[2233] = -288;
    mem[2234] = -289;
    mem[2235] = -291;
    mem[2236] = -292;
    mem[2237] = -294;
    mem[2238] = -295;
    mem[2239] = -297;
    mem[2240] = -298;
    mem[2241] = -300;
    mem[2242] = -301;
    mem[2243] = -303;
    mem[2244] = -304;
    mem[2245] = -306;
    mem[2246] = -307;
    mem[2247] = -309;
    mem[2248] = -310;
    mem[2249] = -312;
    mem[2250] = -313;
    mem[2251] = -315;
    mem[2252] = -316;
    mem[2253] = -318;
    mem[2254] = -319;
    mem[2255] = -321;
    mem[2256] = -322;
    mem[2257] = -324;
    mem[2258] = -325;
    mem[2259] = -327;
    mem[2260] = -328;
    mem[2261] = -329;
    mem[2262] = -331;
    mem[2263] = -332;
    mem[2264] = -334;
    mem[2265] = -335;
    mem[2266] = -337;
    mem[2267] = -338;
    mem[2268] = -340;
    mem[2269] = -341;
    mem[2270] = -343;
    mem[2271] = -344;
    mem[2272] = -346;
    mem[2273] = -347;
    mem[2274] = -349;
    mem[2275] = -350;
    mem[2276] = -352;
    mem[2277] = -353;
    mem[2278] = -355;
    mem[2279] = -356;
    mem[2280] = -358;
    mem[2281] = -359;
    mem[2282] = -361;
    mem[2283] = -362;
    mem[2284] = -363;
    mem[2285] = -365;
    mem[2286] = -366;
    mem[2287] = -368;
    mem[2288] = -369;
    mem[2289] = -371;
    mem[2290] = -372;
    mem[2291] = -374;
    mem[2292] = -375;
    mem[2293] = -377;
    mem[2294] = -378;
    mem[2295] = -380;
    mem[2296] = -381;
    mem[2297] = -383;
    mem[2298] = -384;
    mem[2299] = -385;
    mem[2300] = -387;
    mem[2301] = -388;
    mem[2302] = -390;
    mem[2303] = -391;
    mem[2304] = -393;
    mem[2305] = -394;
    mem[2306] = -396;
    mem[2307] = -397;
    mem[2308] = -398;
    mem[2309] = -400;
    mem[2310] = -401;
    mem[2311] = -403;
    mem[2312] = -404;
    mem[2313] = -406;
    mem[2314] = -407;
    mem[2315] = -409;
    mem[2316] = -410;
    mem[2317] = -411;
    mem[2318] = -413;
    mem[2319] = -414;
    mem[2320] = -416;
    mem[2321] = -417;
    mem[2322] = -419;
    mem[2323] = -420;
    mem[2324] = -422;
    mem[2325] = -423;
    mem[2326] = -424;
    mem[2327] = -426;
    mem[2328] = -427;
    mem[2329] = -429;
    mem[2330] = -430;
    mem[2331] = -432;
    mem[2332] = -433;
    mem[2333] = -434;
    mem[2334] = -436;
    mem[2335] = -437;
    mem[2336] = -439;
    mem[2337] = -440;
    mem[2338] = -441;
    mem[2339] = -443;
    mem[2340] = -444;
    mem[2341] = -446;
    mem[2342] = -447;
    mem[2343] = -449;
    mem[2344] = -450;
    mem[2345] = -451;
    mem[2346] = -453;
    mem[2347] = -454;
    mem[2348] = -456;
    mem[2349] = -457;
    mem[2350] = -458;
    mem[2351] = -460;
    mem[2352] = -461;
    mem[2353] = -463;
    mem[2354] = -464;
    mem[2355] = -465;
    mem[2356] = -467;
    mem[2357] = -468;
    mem[2358] = -470;
    mem[2359] = -471;
    mem[2360] = -472;
    mem[2361] = -474;
    mem[2362] = -475;
    mem[2363] = -477;
    mem[2364] = -478;
    mem[2365] = -479;
    mem[2366] = -481;
    mem[2367] = -482;
    mem[2368] = -484;
    mem[2369] = -485;
    mem[2370] = -486;
    mem[2371] = -488;
    mem[2372] = -489;
    mem[2373] = -490;
    mem[2374] = -492;
    mem[2375] = -493;
    mem[2376] = -495;
    mem[2377] = -496;
    mem[2378] = -497;
    mem[2379] = -499;
    mem[2380] = -500;
    mem[2381] = -501;
    mem[2382] = -503;
    mem[2383] = -504;
    mem[2384] = -506;
    mem[2385] = -507;
    mem[2386] = -508;
    mem[2387] = -510;
    mem[2388] = -511;
    mem[2389] = -512;
    mem[2390] = -514;
    mem[2391] = -515;
    mem[2392] = -516;
    mem[2393] = -518;
    mem[2394] = -519;
    mem[2395] = -520;
    mem[2396] = -522;
    mem[2397] = -523;
    mem[2398] = -525;
    mem[2399] = -526;
    mem[2400] = -527;
    mem[2401] = -529;
    mem[2402] = -530;
    mem[2403] = -531;
    mem[2404] = -533;
    mem[2405] = -534;
    mem[2406] = -535;
    mem[2407] = -537;
    mem[2408] = -538;
    mem[2409] = -539;
    mem[2410] = -541;
    mem[2411] = -542;
    mem[2412] = -543;
    mem[2413] = -545;
    mem[2414] = -546;
    mem[2415] = -547;
    mem[2416] = -549;
    mem[2417] = -550;
    mem[2418] = -551;
    mem[2419] = -553;
    mem[2420] = -554;
    mem[2421] = -555;
    mem[2422] = -557;
    mem[2423] = -558;
    mem[2424] = -559;
    mem[2425] = -561;
    mem[2426] = -562;
    mem[2427] = -563;
    mem[2428] = -564;
    mem[2429] = -566;
    mem[2430] = -567;
    mem[2431] = -568;
    mem[2432] = -570;
    mem[2433] = -571;
    mem[2434] = -572;
    mem[2435] = -574;
    mem[2436] = -575;
    mem[2437] = -576;
    mem[2438] = -577;
    mem[2439] = -579;
    mem[2440] = -580;
    mem[2441] = -581;
    mem[2442] = -583;
    mem[2443] = -584;
    mem[2444] = -585;
    mem[2445] = -587;
    mem[2446] = -588;
    mem[2447] = -589;
    mem[2448] = -590;
    mem[2449] = -592;
    mem[2450] = -593;
    mem[2451] = -594;
    mem[2452] = -596;
    mem[2453] = -597;
    mem[2454] = -598;
    mem[2455] = -599;
    mem[2456] = -601;
    mem[2457] = -602;
    mem[2458] = -603;
    mem[2459] = -604;
    mem[2460] = -606;
    mem[2461] = -607;
    mem[2462] = -608;
    mem[2463] = -609;
    mem[2464] = -611;
    mem[2465] = -612;
    mem[2466] = -613;
    mem[2467] = -615;
    mem[2468] = -616;
    mem[2469] = -617;
    mem[2470] = -618;
    mem[2471] = -620;
    mem[2472] = -621;
    mem[2473] = -622;
    mem[2474] = -623;
    mem[2475] = -625;
    mem[2476] = -626;
    mem[2477] = -627;
    mem[2478] = -628;
    mem[2479] = -630;
    mem[2480] = -631;
    mem[2481] = -632;
    mem[2482] = -633;
    mem[2483] = -634;
    mem[2484] = -636;
    mem[2485] = -637;
    mem[2486] = -638;
    mem[2487] = -639;
    mem[2488] = -641;
    mem[2489] = -642;
    mem[2490] = -643;
    mem[2491] = -644;
    mem[2492] = -645;
    mem[2493] = -647;
    mem[2494] = -648;
    mem[2495] = -649;
    mem[2496] = -650;
    mem[2497] = -652;
    mem[2498] = -653;
    mem[2499] = -654;
    mem[2500] = -655;
    mem[2501] = -656;
    mem[2502] = -658;
    mem[2503] = -659;
    mem[2504] = -660;
    mem[2505] = -661;
    mem[2506] = -662;
    mem[2507] = -664;
    mem[2508] = -665;
    mem[2509] = -666;
    mem[2510] = -667;
    mem[2511] = -668;
    mem[2512] = -670;
    mem[2513] = -671;
    mem[2514] = -672;
    mem[2515] = -673;
    mem[2516] = -674;
    mem[2517] = -676;
    mem[2518] = -677;
    mem[2519] = -678;
    mem[2520] = -679;
    mem[2521] = -680;
    mem[2522] = -681;
    mem[2523] = -683;
    mem[2524] = -684;
    mem[2525] = -685;
    mem[2526] = -686;
    mem[2527] = -687;
    mem[2528] = -688;
    mem[2529] = -690;
    mem[2530] = -691;
    mem[2531] = -692;
    mem[2532] = -693;
    mem[2533] = -694;
    mem[2534] = -695;
    mem[2535] = -696;
    mem[2536] = -698;
    mem[2537] = -699;
    mem[2538] = -700;
    mem[2539] = -701;
    mem[2540] = -702;
    mem[2541] = -703;
    mem[2542] = -705;
    mem[2543] = -706;
    mem[2544] = -707;
    mem[2545] = -708;
    mem[2546] = -709;
    mem[2547] = -710;
    mem[2548] = -711;
    mem[2549] = -712;
    mem[2550] = -714;
    mem[2551] = -715;
    mem[2552] = -716;
    mem[2553] = -717;
    mem[2554] = -718;
    mem[2555] = -719;
    mem[2556] = -720;
    mem[2557] = -721;
    mem[2558] = -723;
    mem[2559] = -724;
    mem[2560] = -725;
    mem[2561] = -726;
    mem[2562] = -727;
    mem[2563] = -728;
    mem[2564] = -729;
    mem[2565] = -730;
    mem[2566] = -731;
    mem[2567] = -732;
    mem[2568] = -734;
    mem[2569] = -735;
    mem[2570] = -736;
    mem[2571] = -737;
    mem[2572] = -738;
    mem[2573] = -739;
    mem[2574] = -740;
    mem[2575] = -741;
    mem[2576] = -742;
    mem[2577] = -743;
    mem[2578] = -744;
    mem[2579] = -746;
    mem[2580] = -747;
    mem[2581] = -748;
    mem[2582] = -749;
    mem[2583] = -750;
    mem[2584] = -751;
    mem[2585] = -752;
    mem[2586] = -753;
    mem[2587] = -754;
    mem[2588] = -755;
    mem[2589] = -756;
    mem[2590] = -757;
    mem[2591] = -758;
    mem[2592] = -759;
    mem[2593] = -760;
    mem[2594] = -762;
    mem[2595] = -763;
    mem[2596] = -764;
    mem[2597] = -765;
    mem[2598] = -766;
    mem[2599] = -767;
    mem[2600] = -768;
    mem[2601] = -769;
    mem[2602] = -770;
    mem[2603] = -771;
    mem[2604] = -772;
    mem[2605] = -773;
    mem[2606] = -774;
    mem[2607] = -775;
    mem[2608] = -776;
    mem[2609] = -777;
    mem[2610] = -778;
    mem[2611] = -779;
    mem[2612] = -780;
    mem[2613] = -781;
    mem[2614] = -782;
    mem[2615] = -783;
    mem[2616] = -784;
    mem[2617] = -785;
    mem[2618] = -786;
    mem[2619] = -787;
    mem[2620] = -788;
    mem[2621] = -789;
    mem[2622] = -790;
    mem[2623] = -791;
    mem[2624] = -792;
    mem[2625] = -793;
    mem[2626] = -794;
    mem[2627] = -795;
    mem[2628] = -796;
    mem[2629] = -797;
    mem[2630] = -798;
    mem[2631] = -799;
    mem[2632] = -800;
    mem[2633] = -801;
    mem[2634] = -802;
    mem[2635] = -803;
    mem[2636] = -804;
    mem[2637] = -805;
    mem[2638] = -806;
    mem[2639] = -807;
    mem[2640] = -808;
    mem[2641] = -809;
    mem[2642] = -810;
    mem[2643] = -811;
    mem[2644] = -812;
    mem[2645] = -813;
    mem[2646] = -814;
    mem[2647] = -815;
    mem[2648] = -816;
    mem[2649] = -817;
    mem[2650] = -817;
    mem[2651] = -818;
    mem[2652] = -819;
    mem[2653] = -820;
    mem[2654] = -821;
    mem[2655] = -822;
    mem[2656] = -823;
    mem[2657] = -824;
    mem[2658] = -825;
    mem[2659] = -826;
    mem[2660] = -827;
    mem[2661] = -828;
    mem[2662] = -829;
    mem[2663] = -830;
    mem[2664] = -831;
    mem[2665] = -831;
    mem[2666] = -832;
    mem[2667] = -833;
    mem[2668] = -834;
    mem[2669] = -835;
    mem[2670] = -836;
    mem[2671] = -837;
    mem[2672] = -838;
    mem[2673] = -839;
    mem[2674] = -840;
    mem[2675] = -840;
    mem[2676] = -841;
    mem[2677] = -842;
    mem[2678] = -843;
    mem[2679] = -844;
    mem[2680] = -845;
    mem[2681] = -846;
    mem[2682] = -847;
    mem[2683] = -848;
    mem[2684] = -848;
    mem[2685] = -849;
    mem[2686] = -850;
    mem[2687] = -851;
    mem[2688] = -852;
    mem[2689] = -853;
    mem[2690] = -854;
    mem[2691] = -855;
    mem[2692] = -855;
    mem[2693] = -856;
    mem[2694] = -857;
    mem[2695] = -858;
    mem[2696] = -859;
    mem[2697] = -860;
    mem[2698] = -861;
    mem[2699] = -861;
    mem[2700] = -862;
    mem[2701] = -863;
    mem[2702] = -864;
    mem[2703] = -865;
    mem[2704] = -866;
    mem[2705] = -867;
    mem[2706] = -867;
    mem[2707] = -868;
    mem[2708] = -869;
    mem[2709] = -870;
    mem[2710] = -871;
    mem[2711] = -872;
    mem[2712] = -872;
    mem[2713] = -873;
    mem[2714] = -874;
    mem[2715] = -875;
    mem[2716] = -876;
    mem[2717] = -876;
    mem[2718] = -877;
    mem[2719] = -878;
    mem[2720] = -879;
    mem[2721] = -880;
    mem[2722] = -880;
    mem[2723] = -881;
    mem[2724] = -882;
    mem[2725] = -883;
    mem[2726] = -884;
    mem[2727] = -884;
    mem[2728] = -885;
    mem[2729] = -886;
    mem[2730] = -887;
    mem[2731] = -888;
    mem[2732] = -888;
    mem[2733] = -889;
    mem[2734] = -890;
    mem[2735] = -891;
    mem[2736] = -891;
    mem[2737] = -892;
    mem[2738] = -893;
    mem[2739] = -894;
    mem[2740] = -895;
    mem[2741] = -895;
    mem[2742] = -896;
    mem[2743] = -897;
    mem[2744] = -898;
    mem[2745] = -898;
    mem[2746] = -899;
    mem[2747] = -900;
    mem[2748] = -901;
    mem[2749] = -901;
    mem[2750] = -902;
    mem[2751] = -903;
    mem[2752] = -904;
    mem[2753] = -904;
    mem[2754] = -905;
    mem[2755] = -906;
    mem[2756] = -907;
    mem[2757] = -907;
    mem[2758] = -908;
    mem[2759] = -909;
    mem[2760] = -909;
    mem[2761] = -910;
    mem[2762] = -911;
    mem[2763] = -912;
    mem[2764] = -912;
    mem[2765] = -913;
    mem[2766] = -914;
    mem[2767] = -914;
    mem[2768] = -915;
    mem[2769] = -916;
    mem[2770] = -917;
    mem[2771] = -917;
    mem[2772] = -918;
    mem[2773] = -919;
    mem[2774] = -919;
    mem[2775] = -920;
    mem[2776] = -921;
    mem[2777] = -921;
    mem[2778] = -922;
    mem[2779] = -923;
    mem[2780] = -923;
    mem[2781] = -924;
    mem[2782] = -925;
    mem[2783] = -925;
    mem[2784] = -926;
    mem[2785] = -927;
    mem[2786] = -927;
    mem[2787] = -928;
    mem[2788] = -929;
    mem[2789] = -929;
    mem[2790] = -930;
    mem[2791] = -931;
    mem[2792] = -931;
    mem[2793] = -932;
    mem[2794] = -933;
    mem[2795] = -933;
    mem[2796] = -934;
    mem[2797] = -935;
    mem[2798] = -935;
    mem[2799] = -936;
    mem[2800] = -937;
    mem[2801] = -937;
    mem[2802] = -938;
    mem[2803] = -938;
    mem[2804] = -939;
    mem[2805] = -940;
    mem[2806] = -940;
    mem[2807] = -941;
    mem[2808] = -942;
    mem[2809] = -942;
    mem[2810] = -943;
    mem[2811] = -943;
    mem[2812] = -944;
    mem[2813] = -945;
    mem[2814] = -945;
    mem[2815] = -946;
    mem[2816] = -946;
    mem[2817] = -947;
    mem[2818] = -948;
    mem[2819] = -948;
    mem[2820] = -949;
    mem[2821] = -949;
    mem[2822] = -950;
    mem[2823] = -951;
    mem[2824] = -951;
    mem[2825] = -952;
    mem[2826] = -952;
    mem[2827] = -953;
    mem[2828] = -954;
    mem[2829] = -954;
    mem[2830] = -955;
    mem[2831] = -955;
    mem[2832] = -956;
    mem[2833] = -956;
    mem[2834] = -957;
    mem[2835] = -957;
    mem[2836] = -958;
    mem[2837] = -959;
    mem[2838] = -959;
    mem[2839] = -960;
    mem[2840] = -960;
    mem[2841] = -961;
    mem[2842] = -961;
    mem[2843] = -962;
    mem[2844] = -962;
    mem[2845] = -963;
    mem[2846] = -963;
    mem[2847] = -964;
    mem[2848] = -965;
    mem[2849] = -965;
    mem[2850] = -966;
    mem[2851] = -966;
    mem[2852] = -967;
    mem[2853] = -967;
    mem[2854] = -968;
    mem[2855] = -968;
    mem[2856] = -969;
    mem[2857] = -969;
    mem[2858] = -970;
    mem[2859] = -970;
    mem[2860] = -971;
    mem[2861] = -971;
    mem[2862] = -972;
    mem[2863] = -972;
    mem[2864] = -973;
    mem[2865] = -973;
    mem[2866] = -974;
    mem[2867] = -974;
    mem[2868] = -975;
    mem[2869] = -975;
    mem[2870] = -976;
    mem[2871] = -976;
    mem[2872] = -977;
    mem[2873] = -977;
    mem[2874] = -977;
    mem[2875] = -978;
    mem[2876] = -978;
    mem[2877] = -979;
    mem[2878] = -979;
    mem[2879] = -980;
    mem[2880] = -980;
    mem[2881] = -981;
    mem[2882] = -981;
    mem[2883] = -982;
    mem[2884] = -982;
    mem[2885] = -982;
    mem[2886] = -983;
    mem[2887] = -983;
    mem[2888] = -984;
    mem[2889] = -984;
    mem[2890] = -985;
    mem[2891] = -985;
    mem[2892] = -986;
    mem[2893] = -986;
    mem[2894] = -986;
    mem[2895] = -987;
    mem[2896] = -987;
    mem[2897] = -988;
    mem[2898] = -988;
    mem[2899] = -988;
    mem[2900] = -989;
    mem[2901] = -989;
    mem[2902] = -990;
    mem[2903] = -990;
    mem[2904] = -990;
    mem[2905] = -991;
    mem[2906] = -991;
    mem[2907] = -992;
    mem[2908] = -992;
    mem[2909] = -992;
    mem[2910] = -993;
    mem[2911] = -993;
    mem[2912] = -994;
    mem[2913] = -994;
    mem[2914] = -994;
    mem[2915] = -995;
    mem[2916] = -995;
    mem[2917] = -995;
    mem[2918] = -996;
    mem[2919] = -996;
    mem[2920] = -997;
    mem[2921] = -997;
    mem[2922] = -997;
    mem[2923] = -998;
    mem[2924] = -998;
    mem[2925] = -998;
    mem[2926] = -999;
    mem[2927] = -999;
    mem[2928] = -999;
    mem[2929] = -1000;
    mem[2930] = -1000;
    mem[2931] = -1000;
    mem[2932] = -1001;
    mem[2933] = -1001;
    mem[2934] = -1001;
    mem[2935] = -1002;
    mem[2936] = -1002;
    mem[2937] = -1002;
    mem[2938] = -1003;
    mem[2939] = -1003;
    mem[2940] = -1003;
    mem[2941] = -1004;
    mem[2942] = -1004;
    mem[2943] = -1004;
    mem[2944] = -1005;
    mem[2945] = -1005;
    mem[2946] = -1005;
    mem[2947] = -1005;
    mem[2948] = -1006;
    mem[2949] = -1006;
    mem[2950] = -1006;
    mem[2951] = -1007;
    mem[2952] = -1007;
    mem[2953] = -1007;
    mem[2954] = -1007;
    mem[2955] = -1008;
    mem[2956] = -1008;
    mem[2957] = -1008;
    mem[2958] = -1009;
    mem[2959] = -1009;
    mem[2960] = -1009;
    mem[2961] = -1009;
    mem[2962] = -1010;
    mem[2963] = -1010;
    mem[2964] = -1010;
    mem[2965] = -1010;
    mem[2966] = -1011;
    mem[2967] = -1011;
    mem[2968] = -1011;
    mem[2969] = -1011;
    mem[2970] = -1012;
    mem[2971] = -1012;
    mem[2972] = -1012;
    mem[2973] = -1012;
    mem[2974] = -1013;
    mem[2975] = -1013;
    mem[2976] = -1013;
    mem[2977] = -1013;
    mem[2978] = -1014;
    mem[2979] = -1014;
    mem[2980] = -1014;
    mem[2981] = -1014;
    mem[2982] = -1014;
    mem[2983] = -1015;
    mem[2984] = -1015;
    mem[2985] = -1015;
    mem[2986] = -1015;
    mem[2987] = -1015;
    mem[2988] = -1016;
    mem[2989] = -1016;
    mem[2990] = -1016;
    mem[2991] = -1016;
    mem[2992] = -1016;
    mem[2993] = -1017;
    mem[2994] = -1017;
    mem[2995] = -1017;
    mem[2996] = -1017;
    mem[2997] = -1017;
    mem[2998] = -1018;
    mem[2999] = -1018;
    mem[3000] = -1018;
    mem[3001] = -1018;
    mem[3002] = -1018;
    mem[3003] = -1018;
    mem[3004] = -1019;
    mem[3005] = -1019;
    mem[3006] = -1019;
    mem[3007] = -1019;
    mem[3008] = -1019;
    mem[3009] = -1019;
    mem[3010] = -1019;
    mem[3011] = -1020;
    mem[3012] = -1020;
    mem[3013] = -1020;
    mem[3014] = -1020;
    mem[3015] = -1020;
    mem[3016] = -1020;
    mem[3017] = -1020;
    mem[3018] = -1021;
    mem[3019] = -1021;
    mem[3020] = -1021;
    mem[3021] = -1021;
    mem[3022] = -1021;
    mem[3023] = -1021;
    mem[3024] = -1021;
    mem[3025] = -1021;
    mem[3026] = -1022;
    mem[3027] = -1022;
    mem[3028] = -1022;
    mem[3029] = -1022;
    mem[3030] = -1022;
    mem[3031] = -1022;
    mem[3032] = -1022;
    mem[3033] = -1022;
    mem[3034] = -1022;
    mem[3035] = -1022;
    mem[3036] = -1023;
    mem[3037] = -1023;
    mem[3038] = -1023;
    mem[3039] = -1023;
    mem[3040] = -1023;
    mem[3041] = -1023;
    mem[3042] = -1023;
    mem[3043] = -1023;
    mem[3044] = -1023;
    mem[3045] = -1023;
    mem[3046] = -1023;
    mem[3047] = -1023;
    mem[3048] = -1023;
    mem[3049] = -1023;
    mem[3050] = -1023;
    mem[3051] = -1024;
    mem[3052] = -1024;
    mem[3053] = -1024;
    mem[3054] = -1024;
    mem[3055] = -1024;
    mem[3056] = -1024;
    mem[3057] = -1024;
    mem[3058] = -1024;
    mem[3059] = -1024;
    mem[3060] = -1024;
    mem[3061] = -1024;
    mem[3062] = -1024;
    mem[3063] = -1024;
    mem[3064] = -1024;
    mem[3065] = -1024;
    mem[3066] = -1024;
    mem[3067] = -1024;
    mem[3068] = -1024;
    mem[3069] = -1024;
    mem[3070] = -1024;
    mem[3071] = -1024;
    mem[3072] = -1024;
    mem[3073] = -1024;
    mem[3074] = -1024;
    mem[3075] = -1024;
    mem[3076] = -1024;
    mem[3077] = -1024;
    mem[3078] = -1024;
    mem[3079] = -1024;
    mem[3080] = -1024;
    mem[3081] = -1024;
    mem[3082] = -1024;
    mem[3083] = -1024;
    mem[3084] = -1024;
    mem[3085] = -1024;
    mem[3086] = -1024;
    mem[3087] = -1024;
    mem[3088] = -1024;
    mem[3089] = -1024;
    mem[3090] = -1024;
    mem[3091] = -1024;
    mem[3092] = -1023;
    mem[3093] = -1023;
    mem[3094] = -1023;
    mem[3095] = -1023;
    mem[3096] = -1023;
    mem[3097] = -1023;
    mem[3098] = -1023;
    mem[3099] = -1023;
    mem[3100] = -1023;
    mem[3101] = -1023;
    mem[3102] = -1023;
    mem[3103] = -1023;
    mem[3104] = -1023;
    mem[3105] = -1023;
    mem[3106] = -1023;
    mem[3107] = -1022;
    mem[3108] = -1022;
    mem[3109] = -1022;
    mem[3110] = -1022;
    mem[3111] = -1022;
    mem[3112] = -1022;
    mem[3113] = -1022;
    mem[3114] = -1022;
    mem[3115] = -1022;
    mem[3116] = -1022;
    mem[3117] = -1021;
    mem[3118] = -1021;
    mem[3119] = -1021;
    mem[3120] = -1021;
    mem[3121] = -1021;
    mem[3122] = -1021;
    mem[3123] = -1021;
    mem[3124] = -1021;
    mem[3125] = -1021;
    mem[3126] = -1020;
    mem[3127] = -1020;
    mem[3128] = -1020;
    mem[3129] = -1020;
    mem[3130] = -1020;
    mem[3131] = -1020;
    mem[3132] = -1020;
    mem[3133] = -1019;
    mem[3134] = -1019;
    mem[3135] = -1019;
    mem[3136] = -1019;
    mem[3137] = -1019;
    mem[3138] = -1019;
    mem[3139] = -1018;
    mem[3140] = -1018;
    mem[3141] = -1018;
    mem[3142] = -1018;
    mem[3143] = -1018;
    mem[3144] = -1018;
    mem[3145] = -1017;
    mem[3146] = -1017;
    mem[3147] = -1017;
    mem[3148] = -1017;
    mem[3149] = -1017;
    mem[3150] = -1017;
    mem[3151] = -1016;
    mem[3152] = -1016;
    mem[3153] = -1016;
    mem[3154] = -1016;
    mem[3155] = -1016;
    mem[3156] = -1015;
    mem[3157] = -1015;
    mem[3158] = -1015;
    mem[3159] = -1015;
    mem[3160] = -1015;
    mem[3161] = -1014;
    mem[3162] = -1014;
    mem[3163] = -1014;
    mem[3164] = -1014;
    mem[3165] = -1013;
    mem[3166] = -1013;
    mem[3167] = -1013;
    mem[3168] = -1013;
    mem[3169] = -1013;
    mem[3170] = -1012;
    mem[3171] = -1012;
    mem[3172] = -1012;
    mem[3173] = -1012;
    mem[3174] = -1011;
    mem[3175] = -1011;
    mem[3176] = -1011;
    mem[3177] = -1011;
    mem[3178] = -1010;
    mem[3179] = -1010;
    mem[3180] = -1010;
    mem[3181] = -1010;
    mem[3182] = -1009;
    mem[3183] = -1009;
    mem[3184] = -1009;
    mem[3185] = -1008;
    mem[3186] = -1008;
    mem[3187] = -1008;
    mem[3188] = -1008;
    mem[3189] = -1007;
    mem[3190] = -1007;
    mem[3191] = -1007;
    mem[3192] = -1006;
    mem[3193] = -1006;
    mem[3194] = -1006;
    mem[3195] = -1006;
    mem[3196] = -1005;
    mem[3197] = -1005;
    mem[3198] = -1005;
    mem[3199] = -1004;
    mem[3200] = -1004;
    mem[3201] = -1004;
    mem[3202] = -1003;
    mem[3203] = -1003;
    mem[3204] = -1003;
    mem[3205] = -1003;
    mem[3206] = -1002;
    mem[3207] = -1002;
    mem[3208] = -1002;
    mem[3209] = -1001;
    mem[3210] = -1001;
    mem[3211] = -1001;
    mem[3212] = -1000;
    mem[3213] = -1000;
    mem[3214] = -1000;
    mem[3215] = -999;
    mem[3216] = -999;
    mem[3217] = -999;
    mem[3218] = -998;
    mem[3219] = -998;
    mem[3220] = -997;
    mem[3221] = -997;
    mem[3222] = -997;
    mem[3223] = -996;
    mem[3224] = -996;
    mem[3225] = -996;
    mem[3226] = -995;
    mem[3227] = -995;
    mem[3228] = -995;
    mem[3229] = -994;
    mem[3230] = -994;
    mem[3231] = -993;
    mem[3232] = -993;
    mem[3233] = -993;
    mem[3234] = -992;
    mem[3235] = -992;
    mem[3236] = -991;
    mem[3237] = -991;
    mem[3238] = -991;
    mem[3239] = -990;
    mem[3240] = -990;
    mem[3241] = -989;
    mem[3242] = -989;
    mem[3243] = -989;
    mem[3244] = -988;
    mem[3245] = -988;
    mem[3246] = -987;
    mem[3247] = -987;
    mem[3248] = -987;
    mem[3249] = -986;
    mem[3250] = -986;
    mem[3251] = -985;
    mem[3252] = -985;
    mem[3253] = -984;
    mem[3254] = -984;
    mem[3255] = -984;
    mem[3256] = -983;
    mem[3257] = -983;
    mem[3258] = -982;
    mem[3259] = -982;
    mem[3260] = -981;
    mem[3261] = -981;
    mem[3262] = -980;
    mem[3263] = -980;
    mem[3264] = -980;
    mem[3265] = -979;
    mem[3266] = -979;
    mem[3267] = -978;
    mem[3268] = -978;
    mem[3269] = -977;
    mem[3270] = -977;
    mem[3271] = -976;
    mem[3272] = -976;
    mem[3273] = -975;
    mem[3274] = -975;
    mem[3275] = -974;
    mem[3276] = -974;
    mem[3277] = -973;
    mem[3278] = -973;
    mem[3279] = -972;
    mem[3280] = -972;
    mem[3281] = -971;
    mem[3282] = -971;
    mem[3283] = -970;
    mem[3284] = -970;
    mem[3285] = -969;
    mem[3286] = -969;
    mem[3287] = -968;
    mem[3288] = -968;
    mem[3289] = -967;
    mem[3290] = -967;
    mem[3291] = -966;
    mem[3292] = -966;
    mem[3293] = -965;
    mem[3294] = -965;
    mem[3295] = -964;
    mem[3296] = -964;
    mem[3297] = -963;
    mem[3298] = -963;
    mem[3299] = -962;
    mem[3300] = -962;
    mem[3301] = -961;
    mem[3302] = -960;
    mem[3303] = -960;
    mem[3304] = -959;
    mem[3305] = -959;
    mem[3306] = -958;
    mem[3307] = -958;
    mem[3308] = -957;
    mem[3309] = -957;
    mem[3310] = -956;
    mem[3311] = -955;
    mem[3312] = -955;
    mem[3313] = -954;
    mem[3314] = -954;
    mem[3315] = -953;
    mem[3316] = -953;
    mem[3317] = -952;
    mem[3318] = -951;
    mem[3319] = -951;
    mem[3320] = -950;
    mem[3321] = -950;
    mem[3322] = -949;
    mem[3323] = -949;
    mem[3324] = -948;
    mem[3325] = -947;
    mem[3326] = -947;
    mem[3327] = -946;
    mem[3328] = -946;
    mem[3329] = -945;
    mem[3330] = -944;
    mem[3331] = -944;
    mem[3332] = -943;
    mem[3333] = -943;
    mem[3334] = -942;
    mem[3335] = -941;
    mem[3336] = -941;
    mem[3337] = -940;
    mem[3338] = -939;
    mem[3339] = -939;
    mem[3340] = -938;
    mem[3341] = -938;
    mem[3342] = -937;
    mem[3343] = -936;
    mem[3344] = -936;
    mem[3345] = -935;
    mem[3346] = -934;
    mem[3347] = -934;
    mem[3348] = -933;
    mem[3349] = -932;
    mem[3350] = -932;
    mem[3351] = -931;
    mem[3352] = -930;
    mem[3353] = -930;
    mem[3354] = -929;
    mem[3355] = -928;
    mem[3356] = -928;
    mem[3357] = -927;
    mem[3358] = -926;
    mem[3359] = -926;
    mem[3360] = -925;
    mem[3361] = -924;
    mem[3362] = -924;
    mem[3363] = -923;
    mem[3364] = -922;
    mem[3365] = -922;
    mem[3366] = -921;
    mem[3367] = -920;
    mem[3368] = -920;
    mem[3369] = -919;
    mem[3370] = -918;
    mem[3371] = -918;
    mem[3372] = -917;
    mem[3373] = -916;
    mem[3374] = -915;
    mem[3375] = -915;
    mem[3376] = -914;
    mem[3377] = -913;
    mem[3378] = -913;
    mem[3379] = -912;
    mem[3380] = -911;
    mem[3381] = -911;
    mem[3382] = -910;
    mem[3383] = -909;
    mem[3384] = -908;
    mem[3385] = -908;
    mem[3386] = -907;
    mem[3387] = -906;
    mem[3388] = -905;
    mem[3389] = -905;
    mem[3390] = -904;
    mem[3391] = -903;
    mem[3392] = -902;
    mem[3393] = -902;
    mem[3394] = -901;
    mem[3395] = -900;
    mem[3396] = -899;
    mem[3397] = -899;
    mem[3398] = -898;
    mem[3399] = -897;
    mem[3400] = -896;
    mem[3401] = -896;
    mem[3402] = -895;
    mem[3403] = -894;
    mem[3404] = -893;
    mem[3405] = -893;
    mem[3406] = -892;
    mem[3407] = -891;
    mem[3408] = -890;
    mem[3409] = -890;
    mem[3410] = -889;
    mem[3411] = -888;
    mem[3412] = -887;
    mem[3413] = -886;
    mem[3414] = -886;
    mem[3415] = -885;
    mem[3416] = -884;
    mem[3417] = -883;
    mem[3418] = -882;
    mem[3419] = -882;
    mem[3420] = -881;
    mem[3421] = -880;
    mem[3422] = -879;
    mem[3423] = -878;
    mem[3424] = -878;
    mem[3425] = -877;
    mem[3426] = -876;
    mem[3427] = -875;
    mem[3428] = -874;
    mem[3429] = -874;
    mem[3430] = -873;
    mem[3431] = -872;
    mem[3432] = -871;
    mem[3433] = -870;
    mem[3434] = -869;
    mem[3435] = -869;
    mem[3436] = -868;
    mem[3437] = -867;
    mem[3438] = -866;
    mem[3439] = -865;
    mem[3440] = -864;
    mem[3441] = -864;
    mem[3442] = -863;
    mem[3443] = -862;
    mem[3444] = -861;
    mem[3445] = -860;
    mem[3446] = -859;
    mem[3447] = -858;
    mem[3448] = -858;
    mem[3449] = -857;
    mem[3450] = -856;
    mem[3451] = -855;
    mem[3452] = -854;
    mem[3453] = -853;
    mem[3454] = -852;
    mem[3455] = -852;
    mem[3456] = -851;
    mem[3457] = -850;
    mem[3458] = -849;
    mem[3459] = -848;
    mem[3460] = -847;
    mem[3461] = -846;
    mem[3462] = -845;
    mem[3463] = -845;
    mem[3464] = -844;
    mem[3465] = -843;
    mem[3466] = -842;
    mem[3467] = -841;
    mem[3468] = -840;
    mem[3469] = -839;
    mem[3470] = -838;
    mem[3471] = -837;
    mem[3472] = -836;
    mem[3473] = -836;
    mem[3474] = -835;
    mem[3475] = -834;
    mem[3476] = -833;
    mem[3477] = -832;
    mem[3478] = -831;
    mem[3479] = -830;
    mem[3480] = -829;
    mem[3481] = -828;
    mem[3482] = -827;
    mem[3483] = -826;
    mem[3484] = -825;
    mem[3485] = -824;
    mem[3486] = -824;
    mem[3487] = -823;
    mem[3488] = -822;
    mem[3489] = -821;
    mem[3490] = -820;
    mem[3491] = -819;
    mem[3492] = -818;
    mem[3493] = -817;
    mem[3494] = -816;
    mem[3495] = -815;
    mem[3496] = -814;
    mem[3497] = -813;
    mem[3498] = -812;
    mem[3499] = -811;
    mem[3500] = -810;
    mem[3501] = -809;
    mem[3502] = -808;
    mem[3503] = -807;
    mem[3504] = -806;
    mem[3505] = -805;
    mem[3506] = -804;
    mem[3507] = -804;
    mem[3508] = -803;
    mem[3509] = -802;
    mem[3510] = -801;
    mem[3511] = -800;
    mem[3512] = -799;
    mem[3513] = -798;
    mem[3514] = -797;
    mem[3515] = -796;
    mem[3516] = -795;
    mem[3517] = -794;
    mem[3518] = -793;
    mem[3519] = -792;
    mem[3520] = -791;
    mem[3521] = -790;
    mem[3522] = -789;
    mem[3523] = -788;
    mem[3524] = -787;
    mem[3525] = -786;
    mem[3526] = -785;
    mem[3527] = -784;
    mem[3528] = -783;
    mem[3529] = -782;
    mem[3530] = -781;
    mem[3531] = -780;
    mem[3532] = -779;
    mem[3533] = -778;
    mem[3534] = -777;
    mem[3535] = -776;
    mem[3536] = -774;
    mem[3537] = -773;
    mem[3538] = -772;
    mem[3539] = -771;
    mem[3540] = -770;
    mem[3541] = -769;
    mem[3542] = -768;
    mem[3543] = -767;
    mem[3544] = -766;
    mem[3545] = -765;
    mem[3546] = -764;
    mem[3547] = -763;
    mem[3548] = -762;
    mem[3549] = -761;
    mem[3550] = -760;
    mem[3551] = -759;
    mem[3552] = -758;
    mem[3553] = -757;
    mem[3554] = -756;
    mem[3555] = -755;
    mem[3556] = -754;
    mem[3557] = -753;
    mem[3558] = -751;
    mem[3559] = -750;
    mem[3560] = -749;
    mem[3561] = -748;
    mem[3562] = -747;
    mem[3563] = -746;
    mem[3564] = -745;
    mem[3565] = -744;
    mem[3566] = -743;
    mem[3567] = -742;
    mem[3568] = -741;
    mem[3569] = -740;
    mem[3570] = -739;
    mem[3571] = -737;
    mem[3572] = -736;
    mem[3573] = -735;
    mem[3574] = -734;
    mem[3575] = -733;
    mem[3576] = -732;
    mem[3577] = -731;
    mem[3578] = -730;
    mem[3579] = -729;
    mem[3580] = -728;
    mem[3581] = -726;
    mem[3582] = -725;
    mem[3583] = -724;
    mem[3584] = -723;
    mem[3585] = -722;
    mem[3586] = -721;
    mem[3587] = -720;
    mem[3588] = -719;
    mem[3589] = -718;
    mem[3590] = -716;
    mem[3591] = -715;
    mem[3592] = -714;
    mem[3593] = -713;
    mem[3594] = -712;
    mem[3595] = -711;
    mem[3596] = -710;
    mem[3597] = -708;
    mem[3598] = -707;
    mem[3599] = -706;
    mem[3600] = -705;
    mem[3601] = -704;
    mem[3602] = -703;
    mem[3603] = -702;
    mem[3604] = -701;
    mem[3605] = -699;
    mem[3606] = -698;
    mem[3607] = -697;
    mem[3608] = -696;
    mem[3609] = -695;
    mem[3610] = -694;
    mem[3611] = -692;
    mem[3612] = -691;
    mem[3613] = -690;
    mem[3614] = -689;
    mem[3615] = -688;
    mem[3616] = -687;
    mem[3617] = -685;
    mem[3618] = -684;
    mem[3619] = -683;
    mem[3620] = -682;
    mem[3621] = -681;
    mem[3622] = -680;
    mem[3623] = -678;
    mem[3624] = -677;
    mem[3625] = -676;
    mem[3626] = -675;
    mem[3627] = -674;
    mem[3628] = -673;
    mem[3629] = -671;
    mem[3630] = -670;
    mem[3631] = -669;
    mem[3632] = -668;
    mem[3633] = -667;
    mem[3634] = -665;
    mem[3635] = -664;
    mem[3636] = -663;
    mem[3637] = -662;
    mem[3638] = -661;
    mem[3639] = -659;
    mem[3640] = -658;
    mem[3641] = -657;
    mem[3642] = -656;
    mem[3643] = -655;
    mem[3644] = -653;
    mem[3645] = -652;
    mem[3646] = -651;
    mem[3647] = -650;
    mem[3648] = -649;
    mem[3649] = -647;
    mem[3650] = -646;
    mem[3651] = -645;
    mem[3652] = -644;
    mem[3653] = -642;
    mem[3654] = -641;
    mem[3655] = -640;
    mem[3656] = -639;
    mem[3657] = -638;
    mem[3658] = -636;
    mem[3659] = -635;
    mem[3660] = -634;
    mem[3661] = -633;
    mem[3662] = -631;
    mem[3663] = -630;
    mem[3664] = -629;
    mem[3665] = -628;
    mem[3666] = -626;
    mem[3667] = -625;
    mem[3668] = -624;
    mem[3669] = -623;
    mem[3670] = -621;
    mem[3671] = -620;
    mem[3672] = -619;
    mem[3673] = -618;
    mem[3674] = -616;
    mem[3675] = -615;
    mem[3676] = -614;
    mem[3677] = -613;
    mem[3678] = -611;
    mem[3679] = -610;
    mem[3680] = -609;
    mem[3681] = -608;
    mem[3682] = -606;
    mem[3683] = -605;
    mem[3684] = -604;
    mem[3685] = -603;
    mem[3686] = -601;
    mem[3687] = -600;
    mem[3688] = -599;
    mem[3689] = -597;
    mem[3690] = -596;
    mem[3691] = -595;
    mem[3692] = -594;
    mem[3693] = -592;
    mem[3694] = -591;
    mem[3695] = -590;
    mem[3696] = -588;
    mem[3697] = -587;
    mem[3698] = -586;
    mem[3699] = -585;
    mem[3700] = -583;
    mem[3701] = -582;
    mem[3702] = -581;
    mem[3703] = -579;
    mem[3704] = -578;
    mem[3705] = -577;
    mem[3706] = -576;
    mem[3707] = -574;
    mem[3708] = -573;
    mem[3709] = -572;
    mem[3710] = -570;
    mem[3711] = -569;
    mem[3712] = -568;
    mem[3713] = -566;
    mem[3714] = -565;
    mem[3715] = -564;
    mem[3716] = -562;
    mem[3717] = -561;
    mem[3718] = -560;
    mem[3719] = -559;
    mem[3720] = -557;
    mem[3721] = -556;
    mem[3722] = -555;
    mem[3723] = -553;
    mem[3724] = -552;
    mem[3725] = -551;
    mem[3726] = -549;
    mem[3727] = -548;
    mem[3728] = -547;
    mem[3729] = -545;
    mem[3730] = -544;
    mem[3731] = -543;
    mem[3732] = -541;
    mem[3733] = -540;
    mem[3734] = -539;
    mem[3735] = -537;
    mem[3736] = -536;
    mem[3737] = -535;
    mem[3738] = -533;
    mem[3739] = -532;
    mem[3740] = -531;
    mem[3741] = -529;
    mem[3742] = -528;
    mem[3743] = -527;
    mem[3744] = -525;
    mem[3745] = -524;
    mem[3746] = -523;
    mem[3747] = -521;
    mem[3748] = -520;
    mem[3749] = -518;
    mem[3750] = -517;
    mem[3751] = -516;
    mem[3752] = -514;
    mem[3753] = -513;
    mem[3754] = -512;
    mem[3755] = -510;
    mem[3756] = -509;
    mem[3757] = -508;
    mem[3758] = -506;
    mem[3759] = -505;
    mem[3760] = -503;
    mem[3761] = -502;
    mem[3762] = -501;
    mem[3763] = -499;
    mem[3764] = -498;
    mem[3765] = -497;
    mem[3766] = -495;
    mem[3767] = -494;
    mem[3768] = -492;
    mem[3769] = -491;
    mem[3770] = -490;
    mem[3771] = -488;
    mem[3772] = -487;
    mem[3773] = -486;
    mem[3774] = -484;
    mem[3775] = -483;
    mem[3776] = -481;
    mem[3777] = -480;
    mem[3778] = -479;
    mem[3779] = -477;
    mem[3780] = -476;
    mem[3781] = -474;
    mem[3782] = -473;
    mem[3783] = -472;
    mem[3784] = -470;
    mem[3785] = -469;
    mem[3786] = -468;
    mem[3787] = -466;
    mem[3788] = -465;
    mem[3789] = -463;
    mem[3790] = -462;
    mem[3791] = -461;
    mem[3792] = -459;
    mem[3793] = -458;
    mem[3794] = -456;
    mem[3795] = -455;
    mem[3796] = -453;
    mem[3797] = -452;
    mem[3798] = -451;
    mem[3799] = -449;
    mem[3800] = -448;
    mem[3801] = -446;
    mem[3802] = -445;
    mem[3803] = -444;
    mem[3804] = -442;
    mem[3805] = -441;
    mem[3806] = -439;
    mem[3807] = -438;
    mem[3808] = -436;
    mem[3809] = -435;
    mem[3810] = -434;
    mem[3811] = -432;
    mem[3812] = -431;
    mem[3813] = -429;
    mem[3814] = -428;
    mem[3815] = -427;
    mem[3816] = -425;
    mem[3817] = -424;
    mem[3818] = -422;
    mem[3819] = -421;
    mem[3820] = -419;
    mem[3821] = -418;
    mem[3822] = -416;
    mem[3823] = -415;
    mem[3824] = -414;
    mem[3825] = -412;
    mem[3826] = -411;
    mem[3827] = -409;
    mem[3828] = -408;
    mem[3829] = -406;
    mem[3830] = -405;
    mem[3831] = -404;
    mem[3832] = -402;
    mem[3833] = -401;
    mem[3834] = -399;
    mem[3835] = -398;
    mem[3836] = -396;
    mem[3837] = -395;
    mem[3838] = -393;
    mem[3839] = -392;
    mem[3840] = -391;
    mem[3841] = -389;
    mem[3842] = -388;
    mem[3843] = -386;
    mem[3844] = -385;
    mem[3845] = -383;
    mem[3846] = -382;
    mem[3847] = -380;
    mem[3848] = -379;
    mem[3849] = -377;
    mem[3850] = -376;
    mem[3851] = -374;
    mem[3852] = -373;
    mem[3853] = -372;
    mem[3854] = -370;
    mem[3855] = -369;
    mem[3856] = -367;
    mem[3857] = -366;
    mem[3858] = -364;
    mem[3859] = -363;
    mem[3860] = -361;
    mem[3861] = -360;
    mem[3862] = -358;
    mem[3863] = -357;
    mem[3864] = -355;
    mem[3865] = -354;
    mem[3866] = -352;
    mem[3867] = -351;
    mem[3868] = -349;
    mem[3869] = -348;
    mem[3870] = -347;
    mem[3871] = -345;
    mem[3872] = -344;
    mem[3873] = -342;
    mem[3874] = -341;
    mem[3875] = -339;
    mem[3876] = -338;
    mem[3877] = -336;
    mem[3878] = -335;
    mem[3879] = -333;
    mem[3880] = -332;
    mem[3881] = -330;
    mem[3882] = -329;
    mem[3883] = -327;
    mem[3884] = -326;
    mem[3885] = -324;
    mem[3886] = -323;
    mem[3887] = -321;
    mem[3888] = -320;
    mem[3889] = -318;
    mem[3890] = -317;
    mem[3891] = -315;
    mem[3892] = -314;
    mem[3893] = -312;
    mem[3894] = -311;
    mem[3895] = -309;
    mem[3896] = -308;
    mem[3897] = -306;
    mem[3898] = -305;
    mem[3899] = -303;
    mem[3900] = -302;
    mem[3901] = -300;
    mem[3902] = -299;
    mem[3903] = -297;
    mem[3904] = -296;
    mem[3905] = -294;
    mem[3906] = -293;
    mem[3907] = -291;
    mem[3908] = -290;
    mem[3909] = -288;
    mem[3910] = -287;
    mem[3911] = -285;
    mem[3912] = -284;
    mem[3913] = -282;
    mem[3914] = -281;
    mem[3915] = -279;
    mem[3916] = -278;
    mem[3917] = -276;
    mem[3918] = -275;
    mem[3919] = -273;
    mem[3920] = -272;
    mem[3921] = -270;
    mem[3922] = -269;
    mem[3923] = -267;
    mem[3924] = -266;
    mem[3925] = -264;
    mem[3926] = -263;
    mem[3927] = -261;
    mem[3928] = -260;
    mem[3929] = -258;
    mem[3930] = -256;
    mem[3931] = -255;
    mem[3932] = -253;
    mem[3933] = -252;
    mem[3934] = -250;
    mem[3935] = -249;
    mem[3936] = -247;
    mem[3937] = -246;
    mem[3938] = -244;
    mem[3939] = -243;
    mem[3940] = -241;
    mem[3941] = -240;
    mem[3942] = -238;
    mem[3943] = -237;
    mem[3944] = -235;
    mem[3945] = -234;
    mem[3946] = -232;
    mem[3947] = -231;
    mem[3948] = -229;
    mem[3949] = -227;
    mem[3950] = -226;
    mem[3951] = -224;
    mem[3952] = -223;
    mem[3953] = -221;
    mem[3954] = -220;
    mem[3955] = -218;
    mem[3956] = -217;
    mem[3957] = -215;
    mem[3958] = -214;
    mem[3959] = -212;
    mem[3960] = -211;
    mem[3961] = -209;
    mem[3962] = -208;
    mem[3963] = -206;
    mem[3964] = -204;
    mem[3965] = -203;
    mem[3966] = -201;
    mem[3967] = -200;
    mem[3968] = -198;
    mem[3969] = -197;
    mem[3970] = -195;
    mem[3971] = -194;
    mem[3972] = -192;
    mem[3973] = -191;
    mem[3974] = -189;
    mem[3975] = -187;
    mem[3976] = -186;
    mem[3977] = -184;
    mem[3978] = -183;
    mem[3979] = -181;
    mem[3980] = -180;
    mem[3981] = -178;
    mem[3982] = -177;
    mem[3983] = -175;
    mem[3984] = -174;
    mem[3985] = -172;
    mem[3986] = -170;
    mem[3987] = -169;
    mem[3988] = -167;
    mem[3989] = -166;
    mem[3990] = -164;
    mem[3991] = -163;
    mem[3992] = -161;
    mem[3993] = -160;
    mem[3994] = -158;
    mem[3995] = -157;
    mem[3996] = -155;
    mem[3997] = -153;
    mem[3998] = -152;
    mem[3999] = -150;
    mem[4000] = -149;
    mem[4001] = -147;
    mem[4002] = -146;
    mem[4003] = -144;
    mem[4004] = -143;
    mem[4005] = -141;
    mem[4006] = -139;
    mem[4007] = -138;
    mem[4008] = -136;
    mem[4009] = -135;
    mem[4010] = -133;
    mem[4011] = -132;
    mem[4012] = -130;
    mem[4013] = -128;
    mem[4014] = -127;
    mem[4015] = -125;
    mem[4016] = -124;
    mem[4017] = -122;
    mem[4018] = -121;
    mem[4019] = -119;
    mem[4020] = -118;
    mem[4021] = -116;
    mem[4022] = -114;
    mem[4023] = -113;
    mem[4024] = -111;
    mem[4025] = -110;
    mem[4026] = -108;
    mem[4027] = -107;
    mem[4028] = -105;
    mem[4029] = -104;
    mem[4030] = -102;
    mem[4031] = -100;
    mem[4032] = -99;
    mem[4033] = -97;
    mem[4034] = -96;
    mem[4035] = -94;
    mem[4036] = -93;
    mem[4037] = -91;
    mem[4038] = -89;
    mem[4039] = -88;
    mem[4040] = -86;
    mem[4041] = -85;
    mem[4042] = -83;
    mem[4043] = -82;
    mem[4044] = -80;
    mem[4045] = -78;
    mem[4046] = -77;
    mem[4047] = -75;
    mem[4048] = -74;
    mem[4049] = -72;
    mem[4050] = -71;
    mem[4051] = -69;
    mem[4052] = -68;
    mem[4053] = -66;
    mem[4054] = -64;
    mem[4055] = -63;
    mem[4056] = -61;
    mem[4057] = -60;
    mem[4058] = -58;
    mem[4059] = -57;
    mem[4060] = -55;
    mem[4061] = -53;
    mem[4062] = -52;
    mem[4063] = -50;
    mem[4064] = -49;
    mem[4065] = -47;
    mem[4066] = -46;
    mem[4067] = -44;
    mem[4068] = -42;
    mem[4069] = -41;
    mem[4070] = -39;
    mem[4071] = -38;
    mem[4072] = -36;
    mem[4073] = -35;
    mem[4074] = -33;
    mem[4075] = -31;
    mem[4076] = -30;
    mem[4077] = -28;
    mem[4078] = -27;
    mem[4079] = -25;
    mem[4080] = -24;
    mem[4081] = -22;
    mem[4082] = -20;
    mem[4083] = -19;
    mem[4084] = -17;
    mem[4085] = -16;
    mem[4086] = -14;
    mem[4087] = -13;
    mem[4088] = -11;
    mem[4089] = -9;
    mem[4090] = -8;
    mem[4091] = -6;
    mem[4092] = -5;
    mem[4093] = -3;
    mem[4094] = -2;
    mem[4095] = 0;
    end
        
    always@(posedge sclk or negedge rst_n)
    if(rst_n == 1'b0)
    data <= 12'b0;
    else if(en == 1'b1)
    data <= mem[addr];
    else 
    data <= 12'b0;
    
endmodule
